module base2log ( // calculo da energia 20 * log10(x) = 6 * log2(x)
    input  logic [31:0] number_i,
    output logic  [7:0] log_o
);
    always @(*) begin
        casex (number_i)
            32'b1???????????????????????????????: log_o = 5'd31 * 6;
            32'b01??????????????????????????????: log_o = 5'd30 * 6;
            32'b001?????????????????????????????: log_o = 5'd29 * 6;
            32'b0001????????????????????????????: log_o = 5'd28 * 6;
            32'b00001???????????????????????????: log_o = 5'd27 * 6;
            32'b000001??????????????????????????: log_o = 5'd26 * 6;
            32'b0000001?????????????????????????: log_o = 5'd25 * 6;
            32'b00000001????????????????????????: log_o = 5'd24 * 6;
            32'b000000001???????????????????????: log_o = 5'd23 * 6;
            32'b0000000001??????????????????????: log_o = 5'd22 * 6;
            32'b00000000001?????????????????????: log_o = 5'd21 * 6;
            32'b000000000001????????????????????: log_o = 5'd20 * 6;
            32'b0000000000001???????????????????: log_o = 5'd19 * 6;
            32'b00000000000001??????????????????: log_o = 5'd18 * 6;
            32'b000000000000001?????????????????: log_o = 5'd17 * 6;
            32'b0000000000000001????????????????: log_o = 5'd16 * 6;
            32'b00000000000000001???????????????: log_o = 5'd15 * 6;
            32'b000000000000000001??????????????: log_o = 5'd14 * 6;
            32'b0000000000000000001?????????????: log_o = 5'd13 * 6;
            32'b00000000000000000001????????????: log_o = 5'd12 * 6;
            32'b000000000000000000001???????????: log_o = 5'd11 * 6;
            32'b0000000000000000000001??????????: log_o = 5'd10 * 6;
            32'b00000000000000000000001?????????: log_o = 5'd9  * 6;
            32'b000000000000000000000001????????: log_o = 5'd8  * 6;
            32'b0000000000000000000000001???????: log_o = 5'd7  * 6;
            32'b00000000000000000000000001??????: log_o = 5'd6  * 6;
            32'b000000000000000000000000001?????: log_o = 5'd5  * 6;
            32'b0000000000000000000000000001????: log_o = 5'd4  * 6;
            32'b00000000000000000000000000001???: log_o = 5'd3  * 6;
            32'b000000000000000000000000000001??: log_o = 5'd2  * 6;
            32'b0000000000000000000000000000001?: log_o = 5'd1  * 6;
            32'b00000000000000000000000000000001: log_o = 5'd0  * 6;
            default: log_o = 5'd0; // zero input
        endcase
    end

endmodule
