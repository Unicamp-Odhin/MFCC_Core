`timescale 1ns/1ps

import mfcc_pkg::mfcc_data_t;

module MFCC_Core #(
    parameter SAMPLE_WIDTH     = 16,       // Largura do sample de áudio
    parameter NUM_COEFFICIENTS = 13,       // Número de coeficientes MFCC
    parameter NUM_FILTERS      = 40,       // Número de filtros Mel
    parameter FRAME_SIZE       = 400,      // Tamanho do quadro de entrada
    parameter FRAME_MOVE       = 160,      // Tamanho do movimento do quadro
    parameter FFT_SIZE         = 512,      // Tamanho da FFT
    parameter PCM_FIFO_DEPTH   = 256,      // Profundidade do FIFO de PCM
    parameter ALPHA            = 16'd31785 // Alpha em Q1.15 (0.97 ≈ 31785)
) (
    input  logic clk,
    input  logic rst_n,

    // audio input
    input  logic [SAMPLE_WIDTH - 1:0] pcm_in,
    input  logic pcm_ready_i,
    
    // control input
    input  logic start_i,

    output logic mfcc_done_o,
    output mfcc_data_t mfcc_data_o [0:NUM_COEFFICIENTS - 1]
);

    logic pre_emphasis_valid;
    logic [SAMPLE_WIDTH - 1:0] pre_emphasized_signal;

    logic fifo_empty, fifo_rd_en;
    logic [SAMPLE_WIDTH - 1:0] fifo_read_data;

    pre_emphasis #(
        .SAMPLE_WIDTH (SAMPLE_WIDTH),
        .ALPHA        (ALPHA) // Alpha em Q1.15 (0.97 ≈ 31785)
    ) u_pre_emphasis (
        .clk          (clk),
        .rst_n        (rst_n),

        .in_valid     (pcm_ready_i),
        .out_valid    (pre_emphasis_valid),

        .x_in         (pcm_in), // Sinal de entrada
        .y_out        (pre_emphasized_signal) // Sinal de saída
    );

    fifo #(
        .DEPTH        (PCM_FIFO_DEPTH),
        .WIDTH        (SAMPLE_WIDTH)
    ) tx_fifo (
        .clk          (clk),
        .rst_n        (rst_n),

        .wr_en_i      (pre_emphasis_valid),
        .rd_en_i      (fifo_rd_en),

        .write_data_i (pre_emphasized_signal),
        .empty_o      (fifo_empty),
        .read_data_o  (fifo_read_data)
    );

    logic [SAMPLE_WIDTH - 1:0] window_buffer_data_o;
    logic window_valid_to_read;
    logic window_rd_en;
    logic start_move;
    logic start_hamming;

    window_buffer #(
        .WIDTH                (SAMPLE_WIDTH),
        .FRAME_SIZE           (FRAME_SIZE),
        .MOVE_SIZE            (FRAME_MOVE)
    ) u_window_buffer (
        .clk                  (clk),                         // 1 bit
        .rst_n                (rst_n),                       // 1 bit

        .start_move           (start_move),                  // 1 bit

        .fifo_rd_en_o         (fifo_rd_en),                  // 1 bit
        .fifo_data_i          (fifo_read_data),              // 16 bits
        .fifo_empty_i         (fifo_empty),                  // 1 bit

        .rd_en_i              (window_rd_en),                // 10 bits
        .read_data_o          (window_buffer_data_o),        // 16 bits
        .valid_to_read_o      (window_valid_to_read),        // 1 bit

        .start_next_state_o   (start_hamming)
    );

    logic hamming_done, hamming_out_valid;
    logic [8:0] frame_ptr;
    logic signed [SAMPLE_WIDTH - 1:0] hamming_sample;

    hamming_window #(
        .SAMPLE_WIDTH     (SAMPLE_WIDTH),
        .NUM_COEFFICIENTS (FRAME_SIZE),
        .NFFT_SIZE        (FFT_SIZE)
    ) u_hamming_window (
        .clk              (clk),
        .rst_n            (rst_n),

        .start_i          (start_hamming),

        .valid_to_read_i  (window_valid_to_read),
        .rd_en_o          (window_rd_en),

        .frame_ptr_o      (frame_ptr),
        .frame_sample_i   (window_buffer_data_o),  // Sinal de entrada
        .hamming_sample_o (hamming_sample),        // Sinal de saída

        .out_valid_o      (hamming_out_valid),
        .done_o           (hamming_done)
    );

    logic [8:0] fft_ptr;
    logic [31:0] fft_power_sample;
    logic fft_power_valid, fft_done;

    fft_radix2 #(
        .NFFT           (FFT_SIZE),
        .INPUT_WIDTH    (SAMPLE_WIDTH),
        .COMPLEX_WIDTH  (SAMPLE_WIDTH * 2)
    ) u_fft (
        .clk            (clk),
        .rst_n          (rst_n),

        .in_valid       (hamming_out_valid),
        .frame_ptr_i    (frame_ptr),
        .real_in        (hamming_sample),

        .start_i        (hamming_done),

        .power_ptr_o    (fft_ptr),
        .power_valid_o  (fft_power_valid),
        .power_sample_o (fft_power_sample),

        .fft_done_o     (fft_done)
    );

    logic mel_done, mel_valid;
    logic [5:0] mel_ptr;
    logic [7:0] mel_sample;

    mel #(
        .NUM_FILTERS                (NUM_FILTERS), 
        .NFFT                       (FFT_SIZE),
        .INPUT_WIDTH                (32),
        .OUTPUT_WIDTH               (8)
    ) u_mel (
        .clk                        (clk),
        .rst_n                      (rst_n),

        .mel_start_i                (fft_done),

        .in_valid                   (fft_power_valid),
        .power_spectrum_frame_ptr   (fft_ptr),
        .power_spectrum_frame_in    (fft_power_sample),

        .mel_done_o                 (mel_done),

        .mel_value_energies         (mel_sample),
        .mel_prt_energies           (mel_ptr),
        .mel_valid                  (mel_valid)
    );

    logic [$clog2(NUM_COEFFICIENTS) - 1:0] ceps_ptr;
    logic [15:0] ceps_sample;
    logic dct_valid, dct_done;
    logic [15:0] coeficientes [0: NUM_COEFFICIENTS - 1];

    dct #(
        .NUM_CEPS    (NUM_COEFFICIENTS),
        .NUM_FILTERS (NUM_FILTERS),
        .INPUT_WIDTH (8),
        .CEPS_WIDTH  (16)
    ) u_dct (
        .clk         (clk),
        .rst_n       (rst_n),

        .in_valid    (mel_valid),
        .frame_ptr_i (mel_ptr),
        .power_in    (mel_sample),
        
        .start_i     (mel_done),

        .dct_done_o  (dct_done),

        .dct_valid_o (dct_valid),
        .ceps_out    (ceps_sample),
        .ceps_ptr_o  (ceps_ptr)
    );

    always_ff @( posedge clk ) begin
        if (dct_valid) begin
            coeficientes[ceps_ptr] <= ceps_sample;
        end
    end

    logic hamming_finished;
    logic idle;
    assign idle = 0;
    //assign idle = (u_window_buffer.current_state == 0); // IDLE state
/*
    always_ff @( posedge clk or negedge rst_n ) begin : RESTARTIG_LOGIC
        if (!rst_n) begin
            start_move       <= 0;
            hamming_finished <= 0;
        end else begin
            if(hamming_done) begin
                hamming_finished <= 1;
            end
            start_move <= hamming_finished && idle;
            if(hamming_finished && idle) begin
                hamming_finished <= 0;
            end
        end
    end
*/

    //assign start_move = hamming_done && idle;
    assign start_move  = start_i;
    //assign start_move  = hamming_done && u_window_buffer.current_state == u_window_buffer.IDLE;
    assign mfcc_done_o = dct_done;
    assign mfcc_data_o = coeficientes;

endmodule
