module MFCC_Core (auto_restart_i,
    clk,
    mfcc_done_o,
    pcm_ready_i,
    rst_n,
    start_i,
    mfcc_data_o,
    pcm_in);
 input auto_restart_i;
 input clk;
 output mfcc_done_o;
 input pcm_ready_i;
 input rst_n;
 input start_i;
 output [207:0] mfcc_data_o;
 input [15:0] pcm_in;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire net2204;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire net2191;
 wire _00577_;
 wire _00578_;
 wire net2190;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire net2189;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire net2187;
 wire net2186;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire net2185;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire net2184;
 wire net2183;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire net2181;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire net2182;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire net2180;
 wire net2179;
 wire _00762_;
 wire net2178;
 wire net2177;
 wire _00765_;
 wire _00766_;
 wire net2176;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire net2171;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire net2170;
 wire net2169;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire net2168;
 wire _01965_;
 wire _01966_;
 wire net2167;
 wire net2172;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire net2166;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire net2164;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire net2163;
 wire _02232_;
 wire net2162;
 wire net2161;
 wire _02235_;
 wire net2160;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire net2158;
 wire _02242_;
 wire net2165;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire net2159;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire net2156;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire net2157;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire net2155;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire net2173;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire net2154;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire net2152;
 wire _02421_;
 wire net2151;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire net2149;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire net2148;
 wire _02444_;
 wire net2147;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire net2146;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire net2145;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire net2144;
 wire _02483_;
 wire net2143;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire net2142;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire net2141;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire net2140;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire net2137;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire net2134;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire net2133;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire net2132;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire net2131;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire net2130;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire net2129;
 wire _03673_;
 wire net2128;
 wire net2126;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire net2125;
 wire _03690_;
 wire _03691_;
 wire net2122;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire net2121;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire net2120;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire net2119;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire net2117;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire net2116;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire net2115;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire net2114;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire net2112;
 wire net2111;
 wire _03871_;
 wire _03872_;
 wire net2110;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire net2109;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire net2106;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire net2104;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire net2103;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire net2105;
 wire _04787_;
 wire _04788_;
 wire net2102;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire net2100;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire net2101;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire net2098;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire net2096;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire net2095;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire net2094;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire net2097;
 wire net2093;
 wire net2092;
 wire net2091;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire net2090;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire net2199;
 wire _05774_;
 wire net2196;
 wire net2195;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire net2194;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire fft_done;
 wire \fft_ptr[0] ;
 wire \fft_ptr[1] ;
 wire \fft_ptr[2] ;
 wire \fft_ptr[3] ;
 wire \fft_ptr[4] ;
 wire \fft_ptr[5] ;
 wire \fft_ptr[6] ;
 wire \fft_ptr[7] ;
 wire \fft_ptr[8] ;
 wire fifo_rd_en;
 wire hamming_done;
 wire hamming_finished;
 wire idle;
 wire mel_done;
 wire \mel_ptr[0] ;
 wire \mel_ptr[1] ;
 wire \mel_ptr[2] ;
 wire \mel_ptr[3] ;
 wire \mel_ptr[4] ;
 wire \mel_ptr[5] ;
 wire mel_valid;
 wire net213;
 wire pre_emphasis_valid;
 wire start_hamming;
 wire start_move;
 wire start_move_auto;
 wire \tx_fifo.read_ptr[0] ;
 wire \tx_fifo.read_ptr[1] ;
 wire \tx_fifo.read_ptr[2] ;
 wire \tx_fifo.read_ptr[3] ;
 wire \tx_fifo.read_ptr[4] ;
 wire \tx_fifo.read_ptr[5] ;
 wire \tx_fifo.read_ptr[6] ;
 wire \tx_fifo.read_ptr[7] ;
 wire \tx_fifo.write_ptr[0] ;
 wire \tx_fifo.write_ptr[1] ;
 wire \tx_fifo.write_ptr[2] ;
 wire \tx_fifo.write_ptr[3] ;
 wire \tx_fifo.write_ptr[4] ;
 wire \tx_fifo.write_ptr[5] ;
 wire \tx_fifo.write_ptr[6] ;
 wire \tx_fifo.write_ptr[7] ;
 wire \u_dct.dct_state[0] ;
 wire \u_dct.dct_state[1] ;
 wire \u_dct.dct_state[2] ;
 wire \u_dct.dct_state[3] ;
 wire \u_dct.k_ptr[0] ;
 wire \u_dct.k_ptr[1] ;
 wire \u_dct.k_ptr[2] ;
 wire \u_dct.k_ptr[3] ;
 wire \u_dct.n_ptr[0] ;
 wire \u_dct.n_ptr[1] ;
 wire \u_dct.n_ptr[2] ;
 wire \u_dct.n_ptr[3] ;
 wire \u_dct.n_ptr[4] ;
 wire \u_dct.n_ptr[5] ;
 wire \u_fft.fft_state[0] ;
 wire \u_fft.fft_state[1] ;
 wire \u_fft.fft_state[2] ;
 wire \u_fft.fft_state[3] ;
 wire \u_fft.power_ptr[0] ;
 wire \u_fft.power_ptr[1] ;
 wire \u_fft.power_ptr[2] ;
 wire \u_fft.power_ptr[3] ;
 wire \u_fft.power_ptr[4] ;
 wire \u_fft.power_ptr[5] ;
 wire \u_fft.power_ptr[6] ;
 wire \u_fft.power_ptr[7] ;
 wire \u_fft.power_ptr[8] ;
 wire \u_fft.power_ptr[9] ;
 wire \u_fft.power_ptr_stage1[0] ;
 wire \u_fft.power_ptr_stage1[1] ;
 wire \u_fft.power_ptr_stage1[2] ;
 wire \u_fft.power_ptr_stage1[3] ;
 wire \u_fft.power_ptr_stage1[4] ;
 wire \u_fft.power_ptr_stage1[5] ;
 wire \u_fft.power_ptr_stage1[6] ;
 wire \u_fft.power_ptr_stage1[7] ;
 wire \u_fft.power_ptr_stage1[8] ;
 wire \u_fft.power_ptr_stage1[9] ;
 wire \u_fft.power_ptr_stage2[0] ;
 wire \u_fft.power_ptr_stage2[1] ;
 wire \u_fft.power_ptr_stage2[2] ;
 wire \u_fft.power_ptr_stage2[3] ;
 wire \u_fft.power_ptr_stage2[4] ;
 wire \u_fft.power_ptr_stage2[5] ;
 wire \u_fft.power_ptr_stage2[6] ;
 wire \u_fft.power_ptr_stage2[7] ;
 wire \u_fft.power_ptr_stage2[8] ;
 wire \u_fft.power_ptr_stage2[9] ;
 wire \u_fft.power_ptr_stage3[0] ;
 wire \u_fft.power_ptr_stage3[1] ;
 wire \u_fft.power_ptr_stage3[2] ;
 wire \u_fft.power_ptr_stage3[3] ;
 wire \u_fft.power_ptr_stage3[4] ;
 wire \u_fft.power_ptr_stage3[5] ;
 wire \u_fft.power_ptr_stage3[6] ;
 wire \u_fft.power_ptr_stage3[7] ;
 wire \u_fft.power_ptr_stage3[8] ;
 wire \u_fft.power_ptr_stage3[9] ;
 wire \u_fft.power_ptr_stage4[9] ;
 wire \u_fft.sched[0] ;
 wire \u_fft.sched[1] ;
 wire \u_fft.sched[20] ;
 wire \u_fft.sched[21] ;
 wire \u_fft.sched[22] ;
 wire \u_fft.sched[23] ;
 wire \u_fft.sched[24] ;
 wire \u_fft.sched[25] ;
 wire \u_fft.sched[26] ;
 wire \u_fft.sched[29] ;
 wire \u_fft.sched[30] ;
 wire \u_fft.sched[31] ;
 wire \u_fft.sched[32] ;
 wire \u_fft.sched[33] ;
 wire \u_fft.sched[34] ;
 wire \u_fft.sched[35] ;
 wire \u_fft.sched[36] ;
 wire \u_fft.sched[37] ;
 wire \u_fft.sched[38] ;
 wire \u_fft.sched[39] ;
 wire \u_fft.sched[40] ;
 wire \u_fft.sched[41] ;
 wire \u_fft.sched[42] ;
 wire \u_fft.sched[43] ;
 wire \u_fft.sched[44] ;
 wire \u_fft.sched[45] ;
 wire \u_fft.sched[46] ;
 wire \u_fft.sched[47] ;
 wire \u_fft.sched[48] ;
 wire \u_fft.sched[49] ;
 wire \u_fft.sched[50] ;
 wire \u_fft.sched[51] ;
 wire \u_fft.sched[52] ;
 wire \u_fft.sched[53] ;
 wire \u_fft.sched[54] ;
 wire \u_fft.sched[55] ;
 wire \u_fft.sched[56] ;
 wire \u_fft.sched[57] ;
 wire \u_fft.sched[58] ;
 wire \u_fft.sched[59] ;
 wire \u_fft.sched[60] ;
 wire \u_fft.sched[61] ;
 wire \u_fft.sched[62] ;
 wire \u_fft.sched[63] ;
 wire \u_fft.sched[64] ;
 wire \u_hamming_window.calc_pointer[0] ;
 wire \u_hamming_window.calc_pointer[10] ;
 wire \u_hamming_window.calc_pointer[11] ;
 wire \u_hamming_window.calc_pointer[12] ;
 wire \u_hamming_window.calc_pointer[13] ;
 wire \u_hamming_window.calc_pointer[14] ;
 wire \u_hamming_window.calc_pointer[15] ;
 wire \u_hamming_window.calc_pointer[16] ;
 wire \u_hamming_window.calc_pointer[17] ;
 wire \u_hamming_window.calc_pointer[18] ;
 wire \u_hamming_window.calc_pointer[19] ;
 wire \u_hamming_window.calc_pointer[1] ;
 wire \u_hamming_window.calc_pointer[20] ;
 wire \u_hamming_window.calc_pointer[21] ;
 wire \u_hamming_window.calc_pointer[22] ;
 wire \u_hamming_window.calc_pointer[23] ;
 wire \u_hamming_window.calc_pointer[24] ;
 wire \u_hamming_window.calc_pointer[25] ;
 wire \u_hamming_window.calc_pointer[26] ;
 wire \u_hamming_window.calc_pointer[27] ;
 wire \u_hamming_window.calc_pointer[28] ;
 wire \u_hamming_window.calc_pointer[29] ;
 wire \u_hamming_window.calc_pointer[2] ;
 wire \u_hamming_window.calc_pointer[30] ;
 wire \u_hamming_window.calc_pointer[31] ;
 wire \u_hamming_window.calc_pointer[3] ;
 wire \u_hamming_window.calc_pointer[4] ;
 wire \u_hamming_window.calc_pointer[5] ;
 wire \u_hamming_window.calc_pointer[6] ;
 wire \u_hamming_window.calc_pointer[7] ;
 wire \u_hamming_window.calc_pointer[8] ;
 wire \u_hamming_window.calc_pointer[9] ;
 wire \u_hamming_window.done ;
 wire \u_hamming_window.frame_ptr[0] ;
 wire \u_hamming_window.frame_ptr[1] ;
 wire \u_hamming_window.frame_ptr[2] ;
 wire \u_hamming_window.frame_ptr[3] ;
 wire \u_hamming_window.frame_ptr[4] ;
 wire \u_hamming_window.frame_ptr[5] ;
 wire \u_hamming_window.frame_ptr[6] ;
 wire \u_hamming_window.frame_ptr[7] ;
 wire \u_hamming_window.frame_ptr[8] ;
 wire \u_hamming_window.hamming_state[0] ;
 wire \u_hamming_window.hamming_state[1] ;
 wire \u_hamming_window.hamming_state[2] ;
 wire \u_hamming_window.hamming_state[3] ;
 wire \u_hamming_window.rd_en_o ;
 wire \u_mel.k[0] ;
 wire \u_mel.k[1] ;
 wire \u_mel.k[2] ;
 wire \u_mel.k[3] ;
 wire \u_mel.k[4] ;
 wire \u_mel.k[5] ;
 wire \u_mel.k[6] ;
 wire \u_mel.k[7] ;
 wire \u_mel.k[8] ;
 wire \u_mel.k_next[0] ;
 wire \u_mel.k_next[1] ;
 wire \u_mel.state[0] ;
 wire \u_mel.state[1] ;
 wire \u_mel.state[2] ;
 wire \u_window_buffer.current_state[0] ;
 wire \u_window_buffer.current_state[2] ;
 wire \u_window_buffer.current_state[3] ;
 wire \u_window_buffer.current_state[4] ;
 wire \u_window_buffer.internal_read_ptr[10] ;
 wire \u_window_buffer.internal_read_ptr[11] ;
 wire \u_window_buffer.internal_read_ptr[12] ;
 wire \u_window_buffer.internal_read_ptr[13] ;
 wire \u_window_buffer.internal_read_ptr[14] ;
 wire \u_window_buffer.internal_read_ptr[15] ;
 wire \u_window_buffer.internal_read_ptr[16] ;
 wire \u_window_buffer.internal_read_ptr[17] ;
 wire \u_window_buffer.internal_read_ptr[18] ;
 wire \u_window_buffer.internal_read_ptr[19] ;
 wire \u_window_buffer.internal_read_ptr[1] ;
 wire \u_window_buffer.internal_read_ptr[20] ;
 wire \u_window_buffer.internal_read_ptr[21] ;
 wire \u_window_buffer.internal_read_ptr[22] ;
 wire \u_window_buffer.internal_read_ptr[23] ;
 wire \u_window_buffer.internal_read_ptr[24] ;
 wire \u_window_buffer.internal_read_ptr[25] ;
 wire \u_window_buffer.internal_read_ptr[26] ;
 wire \u_window_buffer.internal_read_ptr[27] ;
 wire \u_window_buffer.internal_read_ptr[28] ;
 wire \u_window_buffer.internal_read_ptr[29] ;
 wire \u_window_buffer.internal_read_ptr[2] ;
 wire \u_window_buffer.internal_read_ptr[30] ;
 wire \u_window_buffer.internal_read_ptr[31] ;
 wire \u_window_buffer.internal_read_ptr[3] ;
 wire \u_window_buffer.internal_read_ptr[4] ;
 wire \u_window_buffer.internal_read_ptr[5] ;
 wire \u_window_buffer.internal_read_ptr[6] ;
 wire \u_window_buffer.internal_read_ptr[7] ;
 wire \u_window_buffer.internal_read_ptr[8] ;
 wire \u_window_buffer.internal_read_ptr[9] ;
 wire \u_window_buffer.move_counter[0] ;
 wire \u_window_buffer.move_counter[10] ;
 wire \u_window_buffer.move_counter[11] ;
 wire \u_window_buffer.move_counter[12] ;
 wire \u_window_buffer.move_counter[13] ;
 wire \u_window_buffer.move_counter[14] ;
 wire \u_window_buffer.move_counter[15] ;
 wire \u_window_buffer.move_counter[16] ;
 wire \u_window_buffer.move_counter[17] ;
 wire \u_window_buffer.move_counter[18] ;
 wire \u_window_buffer.move_counter[19] ;
 wire \u_window_buffer.move_counter[1] ;
 wire \u_window_buffer.move_counter[20] ;
 wire \u_window_buffer.move_counter[21] ;
 wire \u_window_buffer.move_counter[22] ;
 wire \u_window_buffer.move_counter[23] ;
 wire \u_window_buffer.move_counter[24] ;
 wire \u_window_buffer.move_counter[25] ;
 wire \u_window_buffer.move_counter[26] ;
 wire \u_window_buffer.move_counter[27] ;
 wire \u_window_buffer.move_counter[28] ;
 wire \u_window_buffer.move_counter[29] ;
 wire \u_window_buffer.move_counter[2] ;
 wire \u_window_buffer.move_counter[30] ;
 wire \u_window_buffer.move_counter[31] ;
 wire \u_window_buffer.move_counter[3] ;
 wire \u_window_buffer.move_counter[4] ;
 wire \u_window_buffer.move_counter[5] ;
 wire \u_window_buffer.move_counter[6] ;
 wire \u_window_buffer.move_counter[7] ;
 wire \u_window_buffer.move_counter[8] ;
 wire \u_window_buffer.move_counter[9] ;
 wire \u_window_buffer.next_state_is_valid_to_read ;
 wire \u_window_buffer.read_ptr[0] ;
 wire \u_window_buffer.read_ptr[10] ;
 wire \u_window_buffer.read_ptr[11] ;
 wire \u_window_buffer.read_ptr[12] ;
 wire \u_window_buffer.read_ptr[13] ;
 wire \u_window_buffer.read_ptr[14] ;
 wire \u_window_buffer.read_ptr[15] ;
 wire \u_window_buffer.read_ptr[16] ;
 wire \u_window_buffer.read_ptr[17] ;
 wire \u_window_buffer.read_ptr[18] ;
 wire \u_window_buffer.read_ptr[19] ;
 wire \u_window_buffer.read_ptr[1] ;
 wire \u_window_buffer.read_ptr[20] ;
 wire \u_window_buffer.read_ptr[21] ;
 wire \u_window_buffer.read_ptr[22] ;
 wire \u_window_buffer.read_ptr[23] ;
 wire \u_window_buffer.read_ptr[24] ;
 wire \u_window_buffer.read_ptr[25] ;
 wire \u_window_buffer.read_ptr[26] ;
 wire \u_window_buffer.read_ptr[27] ;
 wire \u_window_buffer.read_ptr[28] ;
 wire \u_window_buffer.read_ptr[29] ;
 wire \u_window_buffer.read_ptr[2] ;
 wire \u_window_buffer.read_ptr[30] ;
 wire \u_window_buffer.read_ptr[31] ;
 wire \u_window_buffer.read_ptr[3] ;
 wire \u_window_buffer.read_ptr[4] ;
 wire \u_window_buffer.read_ptr[5] ;
 wire \u_window_buffer.read_ptr[6] ;
 wire \u_window_buffer.read_ptr[7] ;
 wire \u_window_buffer.read_ptr[8] ;
 wire \u_window_buffer.read_ptr[9] ;
 wire \u_window_buffer.write_ptr[0] ;
 wire \u_window_buffer.write_ptr[10] ;
 wire \u_window_buffer.write_ptr[11] ;
 wire \u_window_buffer.write_ptr[12] ;
 wire \u_window_buffer.write_ptr[13] ;
 wire \u_window_buffer.write_ptr[14] ;
 wire \u_window_buffer.write_ptr[15] ;
 wire \u_window_buffer.write_ptr[16] ;
 wire \u_window_buffer.write_ptr[17] ;
 wire \u_window_buffer.write_ptr[18] ;
 wire \u_window_buffer.write_ptr[19] ;
 wire \u_window_buffer.write_ptr[1] ;
 wire \u_window_buffer.write_ptr[20] ;
 wire \u_window_buffer.write_ptr[21] ;
 wire \u_window_buffer.write_ptr[22] ;
 wire \u_window_buffer.write_ptr[23] ;
 wire \u_window_buffer.write_ptr[24] ;
 wire \u_window_buffer.write_ptr[25] ;
 wire \u_window_buffer.write_ptr[26] ;
 wire \u_window_buffer.write_ptr[27] ;
 wire \u_window_buffer.write_ptr[28] ;
 wire \u_window_buffer.write_ptr[29] ;
 wire \u_window_buffer.write_ptr[2] ;
 wire \u_window_buffer.write_ptr[30] ;
 wire \u_window_buffer.write_ptr[31] ;
 wire \u_window_buffer.write_ptr[3] ;
 wire \u_window_buffer.write_ptr[4] ;
 wire \u_window_buffer.write_ptr[5] ;
 wire \u_window_buffer.write_ptr[6] ;
 wire \u_window_buffer.write_ptr[7] ;
 wire \u_window_buffer.write_ptr[8] ;
 wire \u_window_buffer.write_ptr[9] ;
 wire net2089;
 wire net2099;
 wire net2087;
 wire net2088;
 wire net2084;
 wire net2082;
 wire net2081;
 wire net2078;
 wire net2079;
 wire net2075;
 wire net2073;
 wire net2072;
 wire net2071;
 wire net2069;
 wire net2068;
 wire net2067;
 wire net2066;
 wire net2065;
 wire net2063;
 wire net2062;
 wire net2061;
 wire net2060;
 wire net2059;
 wire net2058;
 wire net2057;
 wire net2056;
 wire net2055;
 wire net2054;
 wire net2053;
 wire net2049;
 wire net2048;
 wire net2047;
 wire net2046;
 wire net2044;
 wire net2043;
 wire net2042;
 wire net2041;
 wire net2040;
 wire net2045;
 wire net2038;
 wire net2037;
 wire net2036;
 wire net2035;
 wire net2034;
 wire net2029;
 wire net2028;
 wire net2026;
 wire net2025;
 wire net2027;
 wire net2024;
 wire net2023;
 wire net2022;
 wire net2021;
 wire net2020;
 wire net2019;
 wire net2018;
 wire net2030;
 wire net2015;
 wire net2014;
 wire net2013;
 wire net2011;
 wire net2010;
 wire net2012;
 wire net2009;
 wire net2008;
 wire net2007;
 wire net2006;
 wire net2005;
 wire net2004;
 wire net2002;
 wire net2001;
 wire net2000;
 wire net1999;
 wire net2003;
 wire net1998;
 wire net1994;
 wire net1993;
 wire net1992;
 wire net1995;
 wire net1990;
 wire net1991;
 wire net1988;
 wire net1984;
 wire net1983;
 wire net1982;
 wire net1981;
 wire net1980;
 wire net1978;
 wire net1977;
 wire net1976;
 wire net1975;
 wire net1973;
 wire net1969;
 wire net1967;
 wire net1965;
 wire net1964;
 wire net1962;
 wire net1963;
 wire net1960;
 wire net1958;
 wire net1957;
 wire net1956;
 wire net1954;
 wire net1952;
 wire net1953;
 wire net1951;
 wire net1950;
 wire net1948;
 wire net1949;
 wire net1947;
 wire net1945;
 wire net1944;
 wire net1943;
 wire net1941;
 wire net1940;
 wire net1939;
 wire net1938;
 wire net1936;
 wire net1934;
 wire net1935;
 wire net1933;
 wire net1932;
 wire net1937;
 wire net1931;
 wire net1930;
 wire net1929;
 wire net1942;
 wire net1928;
 wire net1925;
 wire net1924;
 wire net1923;
 wire net1922;
 wire net1919;
 wire net1917;
 wire net1916;
 wire net1915;
 wire net1914;
 wire net1913;
 wire net1911;
 wire net1908;
 wire net1907;
 wire net1905;
 wire net1903;
 wire net1902;
 wire net1901;
 wire net1904;
 wire net1900;
 wire net1898;
 wire net1906;
 wire net1896;
 wire net1895;
 wire net1894;
 wire net1893;
 wire net1891;
 wire net1892;
 wire net1897;
 wire net1890;
 wire net1889;
 wire net1888;
 wire net1887;
 wire net1886;
 wire net1885;
 wire net1884;
 wire net1883;
 wire net1909;
 wire net1882;
 wire net1880;
 wire net1881;
 wire net1879;
 wire net1877;
 wire net5107;
 wire net1876;
 wire net1875;
 wire net1874;
 wire net1870;
 wire net1871;
 wire net1868;
 wire net5190;
 wire net1864;
 wire net1861;
 wire net1860;
 wire net1859;
 wire net1858;
 wire net1857;
 wire net1856;
 wire net1855;
 wire net1854;
 wire net1850;
 wire net5262;
 wire net1849;
 wire net1848;
 wire net1852;
 wire net1845;
 wire net1844;
 wire net4958;
 wire net1841;
 wire net1840;
 wire net1846;
 wire clknet_leaf_0_clk;
 wire net1842;
 wire net3780;
 wire net3679;
 wire net212;
 wire net211;
 wire net210;
 wire net209;
 wire net5096;
 wire net2198;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2205;
 wire net2206;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2224;
 wire net2226;
 wire net2225;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2236;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2238;
 wire net2240;
 wire net2242;
 wire net2243;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2251;
 wire net2249;
 wire net2250;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2261;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2265;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2266;
 wire net2268;
 wire net2267;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2274;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2296;
 wire net2294;
 wire net2295;
 wire net2297;
 wire net2298;
 wire net2302;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2303;
 wire net2304;
 wire net2310;
 wire net2306;
 wire net2307;
 wire net2309;
 wire net2308;
 wire net2311;
 wire net2312;
 wire net2315;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2322;
 wire net2347;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2327;
 wire net2326;
 wire net2340;
 wire net2328;
 wire net2331;
 wire net2329;
 wire net2330;
 wire net2339;
 wire net2332;
 wire net2335;
 wire net2333;
 wire net2334;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2345;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2346;
 wire net2348;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2356;
 wire net2358;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2375;
 wire net2376;
 wire net2384;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2387;
 wire net2385;
 wire net2386;
 wire net2388;
 wire net2390;
 wire net2389;
 wire net2391;
 wire net2393;
 wire net2396;
 wire net4923;
 wire net2398;
 wire net2397;
 wire net2401;
 wire net2399;
 wire net2400;
 wire net2402;
 wire net2403;
 wire net2409;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2420;
 wire net2412;
 wire net2410;
 wire net2411;
 wire net2413;
 wire net2416;
 wire net2414;
 wire net2415;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2422;
 wire net2421;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2429;
 wire net2430;
 wire net2444;
 wire net2433;
 wire net2432;
 wire net2437;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2438;
 wire net2439;
 wire net2442;
 wire net2440;
 wire net2441;
 wire net2443;
 wire net2445;
 wire net2447;
 wire net2448;
 wire net2450;
 wire net2451;
 wire net2501;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2494;
 wire net2459;
 wire net2483;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2468;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2470;
 wire net2469;
 wire net2471;
 wire net2473;
 wire net2472;
 wire net2475;
 wire net2474;
 wire net2480;
 wire net2476;
 wire net5142;
 wire net2477;
 wire net2479;
 wire net2482;
 wire net2481;
 wire net2484;
 wire net2491;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2492;
 wire net2493;
 wire net2499;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2500;
 wire net2503;
 wire net2507;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2515;
 wire net2516;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2522;
 wire net2521;
 wire net2523;
 wire net2525;
 wire net2524;
 wire net2536;
 wire net2526;
 wire net2527;
 wire net4961;
 wire net2535;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2542;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2543;
 wire net2544;
 wire net2546;
 wire net2547;
 wire net2556;
 wire net2550;
 wire net2548;
 wire net2549;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2557;
 wire net2578;
 wire net2558;
 wire net2577;
 wire net2565;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2570;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2571;
 wire net2576;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2590;
 wire net2589;
 wire net2634;
 wire net2592;
 wire net2593;
 wire net2613;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2609;
 wire net2599;
 wire net2597;
 wire net2598;
 wire net2600;
 wire net2606;
 wire net2605;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2607;
 wire net2608;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2633;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2631;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2630;
 wire net2624;
 wire net2625;
 wire net2627;
 wire net2626;
 wire net2628;
 wire net2629;
 wire net2632;
 wire net2635;
 wire net2637;
 wire net2636;
 wire net2638;
 wire net2644;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2647;
 wire net2645;
 wire net2646;
 wire net2649;
 wire net2648;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2656;
 wire net2664;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2666;
 wire net2667;
 wire net2669;
 wire net2675;
 wire net2674;
 wire net2671;
 wire net2670;
 wire net2672;
 wire net2673;
 wire net2676;
 wire net2678;
 wire net2679;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2691;
 wire net2692;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2712;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2708;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2735;
 wire net2736;
 wire net2738;
 wire net2739;
 wire net2743;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2760;
 wire net2763;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2770;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2782;
 wire net2784;
 wire net2785;
 wire net2787;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2797;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2798;
 wire net2799;
 wire net2802;
 wire net2801;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2809;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2815;
 wire net2816;
 wire net2820;
 wire net2819;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2827;
 wire net2826;
 wire net2828;
 wire net2829;
 wire net2839;
 wire net2832;
 wire net2833;
 wire net2837;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net5089;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2846;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2863;
 wire net2853;
 wire net2854;
 wire net2858;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2869;
 wire net2864;
 wire net2865;
 wire net2868;
 wire net2866;
 wire net2867;
 wire net2870;
 wire net2873;
 wire net2874;
 wire net2877;
 wire net2876;
 wire net2881;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2889;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2897;
 wire net2896;
 wire net2905;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2903;
 wire net2902;
 wire net2904;
 wire net2908;
 wire net2910;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2921;
 wire net2924;
 wire net2923;
 wire net2927;
 wire net2926;
 wire net2929;
 wire net2928;
 wire net2934;
 wire net2930;
 wire net2933;
 wire net2931;
 wire net2932;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2946;
 wire net2947;
 wire net2949;
 wire net2952;
 wire net2950;
 wire net2951;
 wire net2953;
 wire net2954;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2965;
 wire net2986;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2985;
 wire net2975;
 wire net2982;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2983;
 wire net2984;
 wire net2987;
 wire net2988;
 wire net2990;
 wire net2991;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3002;
 wire net3003;
 wire net3005;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3047;
 wire net3037;
 wire net3026;
 wire net3029;
 wire net3027;
 wire net3028;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3050;
 wire net3048;
 wire net3049;
 wire net3051;
 wire net3052;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3090;
 wire net3089;
 wire net3075;
 wire net3068;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3072;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3074;
 wire net3073;
 wire net3083;
 wire net3080;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3081;
 wire net3082;
 wire net3088;
 wire net3084;
 wire net3087;
 wire net3085;
 wire net3086;
 wire net3110;
 wire net3109;
 wire net3091;
 wire net3108;
 wire net3102;
 wire net3093;
 wire net3092;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3107;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3116;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3117;
 wire net3118;
 wire net3123;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3130;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3131;
 wire net3140;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3153;
 wire net3152;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3168;
 wire net3167;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3166;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3169;
 wire net3171;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3186;
 wire net3187;
 wire net3189;
 wire net3190;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3206;
 wire net3204;
 wire net3205;
 wire net3207;
 wire net3224;
 wire net3215;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3214;
 wire net3213;
 wire net3216;
 wire net3217;
 wire net3219;
 wire net3218;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3229;
 wire net3231;
 wire net3230;
 wire net3236;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3237;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3246;
 wire net3248;
 wire net3249;
 wire net3252;
 wire net3250;
 wire net3251;
 wire net3253;
 wire net3259;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3264;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3277;
 wire net3275;
 wire net3276;
 wire net3280;
 wire net3279;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3299;
 wire net3297;
 wire net3298;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3304;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3313;
 wire net3318;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3319;
 wire net3326;
 wire net3323;
 wire net3322;
 wire net3321;
 wire net3324;
 wire net3325;
 wire net3327;
 wire net3328;
 wire net3342;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3340;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3341;
 wire net3343;
 wire net3351;
 wire net3346;
 wire net3345;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3352;
 wire net3353;
 wire net3356;
 wire net3358;
 wire net3359;
 wire net3362;
 wire net3360;
 wire net3361;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3369;
 wire net3377;
 wire net3370;
 wire net3371;
 wire net3375;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3376;
 wire net3378;
 wire net3379;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3387;
 wire net3386;
 wire net3390;
 wire net3395;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3396;
 wire net3397;
 wire net3399;
 wire net3403;
 wire net3405;
 wire net3406;
 wire net3410;
 wire net3411;
 wire net3414;
 wire net3419;
 wire net3420;
 wire net3422;
 wire net3424;
 wire net3444;
 wire net3425;
 wire net3440;
 wire net3426;
 wire net3437;
 wire net3427;
 wire net3428;
 wire net3430;
 wire net3429;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3438;
 wire net3439;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3445;
 wire net3446;
 wire net3452;
 wire net3447;
 wire net3450;
 wire net3448;
 wire net3449;
 wire net3451;
 wire net3457;
 wire net3463;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3464;
 wire net3471;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3479;
 wire net3481;
 wire net3487;
 wire net3488;
 wire net3492;
 wire net3490;
 wire net3491;
 wire net3495;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3509;
 wire net3510;
 wire net3516;
 wire net3512;
 wire net3515;
 wire net3513;
 wire net3514;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3523;
 wire net3528;
 wire net3530;
 wire net3532;
 wire net3535;
 wire net3537;
 wire net3540;
 wire net3541;
 wire net3543;
 wire net3545;
 wire net3547;
 wire net3550;
 wire net3552;
 wire net3554;
 wire net3556;
 wire net3558;
 wire net3560;
 wire net3562;
 wire net3572;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3570;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3571;
 wire net3574;
 wire net3573;
 wire net3575;
 wire net3576;
 wire net3578;
 wire net3579;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3609;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3605;
 wire net3600;
 wire net3599;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3622;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3633;
 wire net3631;
 wire net3632;
 wire net3635;
 wire net3634;
 wire net3640;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3642;
 wire net3641;
 wire net3644;
 wire net3643;
 wire net3647;
 wire net3645;
 wire net3646;
 wire net3648;
 wire net3649;
 wire net3654;
 wire net3652;
 wire net3651;
 wire net3653;
 wire net3657;
 wire net3655;
 wire net3656;
 wire net3660;
 wire net3659;
 wire net3668;
 wire net3661;
 wire net3665;
 wire net3662;
 wire net3663;
 wire net3664;
 wire net3666;
 wire net3667;
 wire net3670;
 wire net3669;
 wire net3672;
 wire net3671;
 wire net3673;
 wire net3674;
 wire net3678;
 wire clknet_leaf_4_clk;
 wire net3680;
 wire clknet_leaf_3_clk;
 wire net3688;
 wire net3681;
 wire net3682;
 wire net3683;
 wire net3686;
 wire net3685;
 wire net3684;
 wire net3687;
 wire clknet_leaf_2_clk;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3694;
 wire net3696;
 wire net3695;
 wire net3698;
 wire net3697;
 wire net3700;
 wire net3699;
 wire net3783;
 wire net3701;
 wire net3702;
 wire net3725;
 wire net3703;
 wire net3704;
 wire net3705;
 wire net3706;
 wire net3707;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3711;
 wire net3712;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3723;
 wire net3724;
 wire net3726;
 wire net3727;
 wire net3728;
 wire net3729;
 wire net3730;
 wire net3731;
 wire net3732;
 wire net3733;
 wire net3782;
 wire net3734;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3781;
 wire net3745;
 wire net3773;
 wire net3746;
 wire net3747;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3753;
 wire net3754;
 wire net3755;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3764;
 wire net3765;
 wire net3766;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3770;
 wire net3771;
 wire net3772;
 wire net3774;
 wire net3775;
 wire net3776;
 wire net3777;
 wire net3778;
 wire net3779;
 wire clknet_leaf_1_clk;
 wire net3784;
 wire net3785;
 wire net1847;
 wire net1853;
 wire net1862;
 wire net1863;
 wire net1866;
 wire net1867;
 wire net1869;
 wire net5203;
 wire net1873;
 wire net1910;
 wire net1912;
 wire net1918;
 wire net1920;
 wire net1921;
 wire net1926;
 wire net1927;
 wire net1946;
 wire net1955;
 wire net1959;
 wire net1961;
 wire net1966;
 wire net1968;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1974;
 wire net1979;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1989;
 wire net1996;
 wire net1997;
 wire net2016;
 wire net2017;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2039;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2064;
 wire net2070;
 wire net2074;
 wire net2076;
 wire net2077;
 wire net2080;
 wire net2083;
 wire net2085;
 wire net2086;
 wire net2107;
 wire net2108;
 wire net2113;
 wire net2118;
 wire net2123;
 wire net2124;
 wire net2127;
 wire net2135;
 wire net2136;
 wire net2138;
 wire net2139;
 wire net2150;
 wire net2153;
 wire net2174;
 wire net2175;
 wire net2188;
 wire net2192;
 wire net2193;
 wire net2207;
 wire net2214;
 wire net2223;
 wire net2230;
 wire net2237;
 wire net2239;
 wire net2241;
 wire net2244;
 wire net2273;
 wire net2275;
 wire net2276;
 wire net2288;
 wire net2305;
 wire net2313;
 wire net2314;
 wire net2316;
 wire net2321;
 wire net2349;
 wire net2350;
 wire net2355;
 wire net2357;
 wire net2359;
 wire net2367;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2377;
 wire net2392;
 wire net2394;
 wire net2428;
 wire net2431;
 wire net2446;
 wire net2449;
 wire net2452;
 wire net2502;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2508;
 wire net2514;
 wire net2517;
 wire net2537;
 wire net2545;
 wire net2582;
 wire net2591;
 wire net2639;
 wire net2650;
 wire net2654;
 wire net2655;
 wire net2665;
 wire net2668;
 wire net2677;
 wire net2680;
 wire net2684;
 wire net2685;
 wire net2690;
 wire net2693;
 wire net2694;
 wire net2722;
 wire net2730;
 wire net2734;
 wire net2737;
 wire net2749;
 wire net2754;
 wire net2759;
 wire net2761;
 wire net2762;
 wire net2764;
 wire net2769;
 wire net2771;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2783;
 wire net2786;
 wire net2788;
 wire net2792;
 wire net2800;
 wire net2808;
 wire net2810;
 wire net2814;
 wire net2817;
 wire net2818;
 wire net2825;
 wire net2830;
 wire net2831;
 wire net2847;
 wire net2871;
 wire net2872;
 wire net2875;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2888;
 wire net2890;
 wire net2891;
 wire net2895;
 wire net2898;
 wire net2906;
 wire net2907;
 wire net2909;
 wire net2911;
 wire net2912;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2922;
 wire net2925;
 wire net2939;
 wire net2944;
 wire net2945;
 wire net2948;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2963;
 wire net2964;
 wire net2966;
 wire net2967;
 wire net2989;
 wire net2992;
 wire net3001;
 wire net3004;
 wire net3006;
 wire net3011;
 wire net3017;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3053;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3132;
 wire net3159;
 wire net3170;
 wire net3172;
 wire net3179;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3188;
 wire net3191;
 wire net3192;
 wire net3228;
 wire net5065;
 wire net3245;
 wire net3247;
 wire net3254;
 wire net3273;
 wire net3274;
 wire net3278;
 wire net3290;
 wire net3296;
 wire net3303;
 wire net3305;
 wire net3306;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3314;
 wire net3320;
 wire net3344;
 wire net3354;
 wire net3355;
 wire net3357;
 wire net3368;
 wire net3380;
 wire net3384;
 wire net3385;
 wire net3388;
 wire net3389;
 wire net3398;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3404;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3412;
 wire net3413;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3421;
 wire net3423;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3458;
 wire net3459;
 wire net3465;
 wire net3478;
 wire net3480;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3489;
 wire net3493;
 wire net3494;
 wire net3496;
 wire net3501;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3511;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3529;
 wire net3531;
 wire net3533;
 wire net3534;
 wire net3536;
 wire net3538;
 wire net3539;
 wire net3542;
 wire net3544;
 wire net3546;
 wire net3548;
 wire net3549;
 wire net3551;
 wire net3553;
 wire net3555;
 wire net3557;
 wire net3559;
 wire net3561;
 wire net3563;
 wire net3577;
 wire net3580;
 wire net3586;
 wire net3613;
 wire net3621;
 wire net3623;
 wire net3627;
 wire net3636;
 wire net3650;
 wire net3658;
 wire net3675;
 wire net3676;
 wire net3677;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net3786;
 wire net3787;
 wire net3788;
 wire net3789;
 wire net3790;
 wire net3791;
 wire net3792;
 wire net3793;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3798;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3832;
 wire net3833;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3841;
 wire net4860;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4864;
 wire net4865;
 wire net4866;
 wire net4867;
 wire net4868;
 wire net4869;
 wire net4870;
 wire net4871;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4888;
 wire net4889;
 wire net4890;
 wire net4891;
 wire net4892;
 wire net4893;
 wire net4894;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4898;
 wire net4899;
 wire net4900;
 wire net4901;
 wire net4902;
 wire net4903;
 wire net4904;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4918;
 wire net4919;
 wire net4920;
 wire net4921;
 wire net4922;
 wire net4924;
 wire net4925;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4932;
 wire net4933;
 wire net4934;
 wire net4962;
 wire net4967;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net5040;
 wire net5041;
 wire net5042;
 wire net5043;
 wire net5044;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5059;
 wire net5060;
 wire net5061;
 wire net5062;
 wire net5063;
 wire net5064;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5069;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5082;
 wire net5083;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5088;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5093;
 wire net5094;
 wire net5095;
 wire net5097;
 wire net5098;
 wire net5099;
 wire net5100;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5111;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5143;
 wire net5144;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5170;
 wire net5171;
 wire net5172;
 wire net5173;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5199;

 sky130_fd_sc_hs__buf_1 place2199 (.A(_04553_),
    .X(net2199));
 sky130_fd_sc_hs__inv_8 _05869_ (.A(net3784),
    .Y(_05774_));
 sky130_fd_sc_hs__buf_1 place2196 (.A(net2195),
    .X(net2196));
 sky130_fd_sc_hs__buf_2 place2195 (.A(_01709_),
    .X(net2195));
 sky130_fd_sc_hs__buf_1 place2204 (.A(_03418_),
    .X(net2204));
 sky130_fd_sc_hs__nor2_1 _05873_ (.A(\u_fft.sched[26] ),
    .B(\u_fft.sched[1] ),
    .Y(_05777_));
 sky130_fd_sc_hs__inv_2 _05874_ (.A(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hs__nor2_1 _05875_ (.A(\u_fft.sched[22] ),
    .B(\u_fft.sched[21] ),
    .Y(_05779_));
 sky130_fd_sc_hs__inv_1 _05876_ (.A(\u_fft.sched[24] ),
    .Y(_05780_));
 sky130_fd_sc_hs__inv_1 _05877_ (.A(\u_fft.sched[23] ),
    .Y(_05781_));
 sky130_fd_sc_hs__inv_2 _05878_ (.A(\u_fft.sched[20] ),
    .Y(_00053_));
 sky130_fd_sc_hs__nand4_1 _05879_ (.A(_05779_),
    .B(_05780_),
    .C(_05781_),
    .D(_00053_),
    .Y(_05782_));
 sky130_fd_sc_hs__nor4_1 _05880_ (.A(\u_fft.sched[0] ),
    .B(\u_fft.sched[25] ),
    .C(_05778_),
    .D(_05782_),
    .Y(_05783_));
 sky130_fd_sc_hs__xnor2_1 _05881_ (.A(\u_fft.sched[29] ),
    .B(_05783_),
    .Y(_00029_));
 sky130_fd_sc_hs__nor3b_1 _05882_ (.A(\u_fft.sched[22] ),
    .B(\u_fft.sched[23] ),
    .C_N(_00055_),
    .Y(_05784_));
 sky130_fd_sc_hs__nor2_1 _05883_ (.A(\u_fft.sched[24] ),
    .B(\u_fft.sched[25] ),
    .Y(_05785_));
 sky130_fd_sc_hs__nand2_1 _05884_ (.A(_05784_),
    .B(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hs__nor2_1 _05885_ (.A(_05778_),
    .B(_05786_),
    .Y(_05787_));
 sky130_fd_sc_hs__xnor2_1 _05886_ (.A(\u_fft.sched[0] ),
    .B(_05787_),
    .Y(_00032_));
 sky130_fd_sc_hs__nor3_1 _05887_ (.A(\u_fft.sched[26] ),
    .B(\u_fft.sched[25] ),
    .C(_05782_),
    .Y(_05788_));
 sky130_fd_sc_hs__xnor2_1 _05888_ (.A(\u_fft.sched[1] ),
    .B(_05788_),
    .Y(_00035_));
 sky130_fd_sc_hs__xor2_1 _05889_ (.A(\u_fft.sched[26] ),
    .B(_05786_),
    .X(_00038_));
 sky130_fd_sc_hs__xor2_1 _05890_ (.A(\u_fft.sched[25] ),
    .B(_05782_),
    .X(_00041_));
 sky130_fd_sc_hs__xnor2_1 _05891_ (.A(\u_fft.sched[24] ),
    .B(_05784_),
    .Y(_00044_));
 sky130_fd_sc_hs__nand2_1 _05892_ (.A(_05779_),
    .B(_00053_),
    .Y(_05789_));
 sky130_fd_sc_hs__xnor2_1 _05893_ (.A(_05781_),
    .B(_05789_),
    .Y(_00047_));
 sky130_fd_sc_hs__xnor2_1 _05894_ (.A(\u_fft.sched[22] ),
    .B(_00055_),
    .Y(_00050_));
 sky130_fd_sc_hs__inv_2 _05895_ (.A(\u_fft.sched[30] ),
    .Y(_00082_));
 sky130_fd_sc_hs__inv_1 _05896_ (.A(\u_fft.sched[31] ),
    .Y(_00083_));
 sky130_fd_sc_hs__nand3b_1 _05897_ (.A_N(\u_fft.sched[32] ),
    .B(_00083_),
    .C(_00082_),
    .Y(_05790_));
 sky130_fd_sc_hs__nor3_1 _05898_ (.A(\u_fft.sched[34] ),
    .B(\u_fft.sched[33] ),
    .C(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hs__inv_1 _05899_ (.A(_05791_),
    .Y(_05792_));
 sky130_fd_sc_hs__nor3_1 _05900_ (.A(\u_fft.sched[36] ),
    .B(\u_fft.sched[35] ),
    .C(_05792_),
    .Y(_05793_));
 sky130_fd_sc_hs__inv_1 _05901_ (.A(\u_fft.sched[38] ),
    .Y(_05794_));
 sky130_fd_sc_hs__inv_1 _05902_ (.A(\u_fft.sched[37] ),
    .Y(_05795_));
 sky130_fd_sc_hs__nand3_1 _05903_ (.A(_05793_),
    .B(_05794_),
    .C(_05795_),
    .Y(_05796_));
 sky130_fd_sc_hs__xor2_1 _05904_ (.A(\u_fft.sched[39] ),
    .B(_05796_),
    .X(_00058_));
 sky130_fd_sc_hs__nor2_1 _05905_ (.A(\u_fft.sched[33] ),
    .B(\u_fft.sched[32] ),
    .Y(_05797_));
 sky130_fd_sc_hs__nand2_1 _05906_ (.A(_05797_),
    .B(_00084_),
    .Y(_05798_));
 sky130_fd_sc_hs__or3_1 _05907_ (.A(\u_fft.sched[35] ),
    .B(\u_fft.sched[34] ),
    .C(_05798_),
    .X(_05799_));
 sky130_fd_sc_hs__nor3_1 _05908_ (.A(\u_fft.sched[37] ),
    .B(\u_fft.sched[36] ),
    .C(_05799_),
    .Y(_05800_));
 sky130_fd_sc_hs__xnor2_1 _05909_ (.A(_05794_),
    .B(_05800_),
    .Y(_00061_));
 sky130_fd_sc_hs__xnor2_1 _05910_ (.A(_05795_),
    .B(_05793_),
    .Y(_00064_));
 sky130_fd_sc_hs__xnor2_1 _05911_ (.A(\u_fft.sched[36] ),
    .B(_05799_),
    .Y(_00067_));
 sky130_fd_sc_hs__xnor2_1 _05912_ (.A(\u_fft.sched[35] ),
    .B(_05792_),
    .Y(_00070_));
 sky130_fd_sc_hs__xnor2_1 _05913_ (.A(\u_fft.sched[34] ),
    .B(_05798_),
    .Y(_00073_));
 sky130_fd_sc_hs__xnor2_1 _05914_ (.A(\u_fft.sched[33] ),
    .B(_05790_),
    .Y(_00076_));
 sky130_fd_sc_hs__xor2_1 _05915_ (.A(\u_fft.sched[32] ),
    .B(_00084_),
    .X(_00079_));
 sky130_fd_sc_hs__clkinv_1 _05916_ (.A(\mel_ptr[3] ),
    .Y(_05801_));
 sky130_fd_sc_hs__inv_1 _05917_ (.A(\mel_ptr[4] ),
    .Y(_05802_));
 sky130_fd_sc_hs__inv_1 _05918_ (.A(\mel_ptr[5] ),
    .Y(_05803_));
 sky130_fd_sc_hs__a21oi_1 _05919_ (.A1(_05801_),
    .A2(_05802_),
    .B1(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hs__buf_4 place2194 (.A(_03427_),
    .X(net2194));
 sky130_fd_sc_hs__nand2_1 _05921_ (.A(net211),
    .B(\u_mel.state[2] ),
    .Y(_05806_));
 sky130_fd_sc_hs__nor2_1 _05922_ (.A(\u_mel.k[3] ),
    .B(\u_mel.k[2] ),
    .Y(_05807_));
 sky130_fd_sc_hs__clkinv_1 _05923_ (.A(\u_mel.k[5] ),
    .Y(_05808_));
 sky130_fd_sc_hs__clkinv_1 _05924_ (.A(\u_mel.k[4] ),
    .Y(_05809_));
 sky130_fd_sc_hs__nand3_1 _05925_ (.A(_05807_),
    .B(_05808_),
    .C(_05809_),
    .Y(_05810_));
 sky130_fd_sc_hs__inv_1 _05926_ (.A(\u_mel.k[7] ),
    .Y(_05811_));
 sky130_fd_sc_hs__inv_1 _05927_ (.A(\u_mel.k[6] ),
    .Y(_05812_));
 sky130_fd_sc_hs__inv_1 _05928_ (.A(\u_mel.k[8] ),
    .Y(_05813_));
 sky130_fd_sc_hs__nand4_1 _05929_ (.A(_05811_),
    .B(_05812_),
    .C(_05813_),
    .D(_00241_),
    .Y(_05814_));
 sky130_fd_sc_hs__nor2_1 _05930_ (.A(_05810_),
    .B(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hs__inv_1 _05931_ (.A(_05815_),
    .Y(_05816_));
 sky130_fd_sc_hs__nor3_1 _05932_ (.A(\mel_ptr[4] ),
    .B(_05801_),
    .C(_05803_),
    .Y(_05817_));
 sky130_fd_sc_hs__inv_1 _05933_ (.A(\mel_ptr[2] ),
    .Y(_05818_));
 sky130_fd_sc_hs__nand3_1 _05934_ (.A(_05817_),
    .B(_05818_),
    .C(_00207_),
    .Y(_05819_));
 sky130_fd_sc_hs__nand2_1 _05935_ (.A(_05819_),
    .B(net211),
    .Y(_05820_));
 sky130_fd_sc_hs__inv_1 _05936_ (.A(_05820_),
    .Y(_05821_));
 sky130_fd_sc_hs__nand2_1 _05937_ (.A(_05821_),
    .B(\u_mel.state[1] ),
    .Y(_05822_));
 sky130_fd_sc_hs__o22ai_1 _05938_ (.A1(_05804_),
    .A2(_05806_),
    .B1(_05816_),
    .B2(_05822_),
    .Y(_00016_));
 sky130_fd_sc_hs__inv_1 _05939_ (.A(\u_mel.state[0] ),
    .Y(_05823_));
 sky130_fd_sc_hs__nand2_1 _05940_ (.A(_05804_),
    .B(\u_mel.state[2] ),
    .Y(_05824_));
 sky130_fd_sc_hs__o211ai_1 _05941_ (.A1(fft_done),
    .A2(_05823_),
    .B1(_05824_),
    .C1(_05821_),
    .Y(_00015_));
 sky130_fd_sc_hs__inv_2 _05942_ (.A(_00237_),
    .Y(_05825_));
 sky130_fd_sc_hs__nor2_1 _05943_ (.A(\u_hamming_window.calc_pointer[6] ),
    .B(\u_hamming_window.calc_pointer[9] ),
    .Y(_05826_));
 sky130_fd_sc_hs__nand3_1 _05944_ (.A(_05826_),
    .B(\u_hamming_window.calc_pointer[4] ),
    .C(\u_hamming_window.calc_pointer[7] ),
    .Y(_05827_));
 sky130_fd_sc_hs__inv_1 _05945_ (.A(\u_hamming_window.calc_pointer[13] ),
    .Y(_05828_));
 sky130_fd_sc_hs__nand2_1 _05946_ (.A(_05828_),
    .B(\u_hamming_window.calc_pointer[8] ),
    .Y(_05829_));
 sky130_fd_sc_hs__inv_2 _05947_ (.A(\u_hamming_window.calc_pointer[15] ),
    .Y(_05830_));
 sky130_fd_sc_hs__inv_1 _05948_ (.A(\u_hamming_window.calc_pointer[14] ),
    .Y(_05831_));
 sky130_fd_sc_hs__nand2_1 _05949_ (.A(_05830_),
    .B(_05831_),
    .Y(_05832_));
 sky130_fd_sc_hs__nor4_1 _05950_ (.A(\u_hamming_window.calc_pointer[12] ),
    .B(\u_hamming_window.calc_pointer[17] ),
    .C(_05829_),
    .D(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hs__inv_2 _05951_ (.A(\u_hamming_window.calc_pointer[2] ),
    .Y(_05834_));
 sky130_fd_sc_hs__inv_1 _05952_ (.A(\u_hamming_window.calc_pointer[5] ),
    .Y(_05835_));
 sky130_fd_sc_hs__nor2_1 _05953_ (.A(\u_hamming_window.calc_pointer[11] ),
    .B(\u_hamming_window.calc_pointer[10] ),
    .Y(_05836_));
 sky130_fd_sc_hs__nand4_1 _05954_ (.A(_05833_),
    .B(_05834_),
    .C(_05835_),
    .D(_05836_),
    .Y(_05837_));
 sky130_fd_sc_hs__nor4_1 _05955_ (.A(\u_hamming_window.calc_pointer[3] ),
    .B(_05825_),
    .C(_05827_),
    .D(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hs__inv_1 _05956_ (.A(\u_hamming_window.calc_pointer[21] ),
    .Y(_05839_));
 sky130_fd_sc_hs__inv_2 _05957_ (.A(\u_hamming_window.calc_pointer[27] ),
    .Y(_05840_));
 sky130_fd_sc_hs__inv_1 _05958_ (.A(\u_hamming_window.calc_pointer[26] ),
    .Y(_05841_));
 sky130_fd_sc_hs__nand2_1 _05959_ (.A(_05840_),
    .B(_05841_),
    .Y(_05842_));
 sky130_fd_sc_hs__inv_2 _05960_ (.A(\u_hamming_window.calc_pointer[24] ),
    .Y(_05843_));
 sky130_fd_sc_hs__inv_1 _05961_ (.A(\u_hamming_window.calc_pointer[29] ),
    .Y(_05844_));
 sky130_fd_sc_hs__inv_2 _05962_ (.A(\u_hamming_window.calc_pointer[28] ),
    .Y(_05845_));
 sky130_fd_sc_hs__inv_1 _05963_ (.A(\u_hamming_window.calc_pointer[30] ),
    .Y(_05846_));
 sky130_fd_sc_hs__nand4_1 _05964_ (.A(_05843_),
    .B(_05844_),
    .C(_05845_),
    .D(_05846_),
    .Y(_05847_));
 sky130_fd_sc_hs__nor3_1 _05965_ (.A(\u_hamming_window.calc_pointer[31] ),
    .B(_05842_),
    .C(_05847_),
    .Y(_05848_));
 sky130_fd_sc_hs__nor2_1 _05966_ (.A(\u_hamming_window.calc_pointer[19] ),
    .B(\u_hamming_window.calc_pointer[18] ),
    .Y(_05849_));
 sky130_fd_sc_hs__inv_2 _05967_ (.A(_05849_),
    .Y(_05850_));
 sky130_fd_sc_hs__clkinv_1 _05968_ (.A(\u_hamming_window.calc_pointer[20] ),
    .Y(_00558_));
 sky130_fd_sc_hs__clkinv_1 _05969_ (.A(\u_hamming_window.calc_pointer[23] ),
    .Y(_00559_));
 sky130_fd_sc_hs__clkinv_1 _05970_ (.A(\u_hamming_window.calc_pointer[22] ),
    .Y(_00560_));
 sky130_fd_sc_hs__clkinv_1 _05971_ (.A(\u_hamming_window.calc_pointer[25] ),
    .Y(_00561_));
 sky130_fd_sc_hs__nand4_1 _05972_ (.A(_00558_),
    .B(_00559_),
    .C(_00560_),
    .D(_00561_),
    .Y(_00562_));
 sky130_fd_sc_hs__nor3_1 _05973_ (.A(\u_hamming_window.calc_pointer[16] ),
    .B(_05850_),
    .C(_00562_),
    .Y(_00563_));
 sky130_fd_sc_hs__nand4_1 _05974_ (.A(_05838_),
    .B(_05839_),
    .C(_05848_),
    .D(_00563_),
    .Y(_00564_));
 sky130_fd_sc_hs__inv_1 _05975_ (.A(\u_hamming_window.hamming_state[0] ),
    .Y(_00565_));
 sky130_fd_sc_hs__inv_1 _05976_ (.A(start_hamming),
    .Y(_00566_));
 sky130_fd_sc_hs__nor2_1 _05977_ (.A(_00565_),
    .B(_00566_),
    .Y(_00567_));
 sky130_fd_sc_hs__a21oi_1 _05978_ (.A1(_00564_),
    .A2(\u_hamming_window.hamming_state[2] ),
    .B1(_00567_),
    .Y(_00568_));
 sky130_fd_sc_hs__nor2_1 _05979_ (.A(net3782),
    .B(_00568_),
    .Y(_00014_));
 sky130_fd_sc_hs__inv_2 _05980_ (.A(\u_dct.n_ptr[3] ),
    .Y(_00569_));
 sky130_fd_sc_hs__nor3_1 _05981_ (.A(\u_dct.n_ptr[2] ),
    .B(\u_dct.n_ptr[4] ),
    .C(_00569_),
    .Y(_00570_));
 sky130_fd_sc_hs__nand3_1 _05982_ (.A(_00570_),
    .B(_00166_),
    .C(\u_dct.n_ptr[5] ),
    .Y(_00571_));
 sky130_fd_sc_hs__nand2_1 _05983_ (.A(_00571_),
    .B(\u_dct.dct_state[2] ),
    .Y(_00572_));
 sky130_fd_sc_hs__nand3_1 _05984_ (.A(\u_dct.k_ptr[2] ),
    .B(\u_dct.k_ptr[3] ),
    .C(_00161_),
    .Y(_00573_));
 sky130_fd_sc_hs__nand2_1 _05985_ (.A(_00573_),
    .B(\u_dct.dct_state[1] ),
    .Y(_00574_));
 sky130_fd_sc_hs__nand2_1 _05986_ (.A(mel_done),
    .B(\u_dct.dct_state[0] ),
    .Y(_00575_));
 sky130_fd_sc_hs__buf_2 place2191 (.A(_05446_),
    .X(net2191));
 sky130_fd_sc_hs__a31oi_1 _05988_ (.A1(_00572_),
    .A2(_00574_),
    .A3(_00575_),
    .B1(net3781),
    .Y(_00008_));
 sky130_fd_sc_hs__inv_2 _05989_ (.A(\u_dct.dct_state[0] ),
    .Y(_00577_));
 sky130_fd_sc_hs__nor2_1 _05990_ (.A(mel_done),
    .B(_00577_),
    .Y(_00578_));
 sky130_fd_sc_hs__buf_1 place2190 (.A(_01689_),
    .X(net2190));
 sky130_fd_sc_hs__inv_2 _05992_ (.A(\u_dct.dct_state[3] ),
    .Y(_00580_));
 sky130_fd_sc_hs__nand3b_1 _05993_ (.A_N(_00578_),
    .B(net211),
    .C(_00580_),
    .Y(_00007_));
 sky130_fd_sc_hs__nand2_1 _05994_ (.A(\u_hamming_window.frame_ptr[7] ),
    .B(\u_hamming_window.frame_ptr[6] ),
    .Y(_00581_));
 sky130_fd_sc_hs__inv_4 _05995_ (.A(\u_hamming_window.frame_ptr[5] ),
    .Y(_00582_));
 sky130_fd_sc_hs__inv_1 _05996_ (.A(\u_hamming_window.frame_ptr[4] ),
    .Y(_00583_));
 sky130_fd_sc_hs__nand2_1 _05997_ (.A(\u_hamming_window.frame_ptr[2] ),
    .B(\u_hamming_window.frame_ptr[1] ),
    .Y(_00584_));
 sky130_fd_sc_hs__nor3b_1 _05998_ (.A(_00583_),
    .B(_00584_),
    .C_N(\u_hamming_window.frame_ptr[3] ),
    .Y(_00585_));
 sky130_fd_sc_hs__nand2_1 _05999_ (.A(_00585_),
    .B(\u_hamming_window.frame_ptr[0] ),
    .Y(_00586_));
 sky130_fd_sc_hs__nor2_1 _06000_ (.A(_00582_),
    .B(_00586_),
    .Y(_00587_));
 sky130_fd_sc_hs__nand3b_1 _06001_ (.A_N(_00581_),
    .B(_00587_),
    .C(\u_hamming_window.frame_ptr[8] ),
    .Y(_00588_));
 sky130_fd_sc_hs__inv_2 _06002_ (.A(\u_hamming_window.hamming_state[2] ),
    .Y(_00589_));
 sky130_fd_sc_hs__nor2_1 _06003_ (.A(_00589_),
    .B(_00564_),
    .Y(_00590_));
 sky130_fd_sc_hs__a21oi_1 _06004_ (.A1(\u_hamming_window.hamming_state[1] ),
    .A2(_00588_),
    .B1(_00590_),
    .Y(_00591_));
 sky130_fd_sc_hs__nor2_1 _06005_ (.A(net3782),
    .B(_00591_),
    .Y(_00013_));
 sky130_fd_sc_hs__inv_2 _06006_ (.A(idle),
    .Y(_00592_));
 sky130_fd_sc_hs__inv_1 _06007_ (.A(start_move),
    .Y(_00593_));
 sky130_fd_sc_hs__nor3_1 _06008_ (.A(_05774_),
    .B(_00592_),
    .C(_00593_),
    .Y(_00006_));
 sky130_fd_sc_hs__buf_1 place2189 (.A(_01713_),
    .X(net2189));
 sky130_fd_sc_hs__xnor2_1 _06010_ (.A(\tx_fifo.write_ptr[4] ),
    .B(\tx_fifo.read_ptr[4] ),
    .Y(_00595_));
 sky130_fd_sc_hs__xnor2_1 _06011_ (.A(\tx_fifo.write_ptr[5] ),
    .B(\tx_fifo.read_ptr[5] ),
    .Y(_00596_));
 sky130_fd_sc_hs__nand2_1 _06012_ (.A(_00595_),
    .B(_00596_),
    .Y(_00597_));
 sky130_fd_sc_hs__inv_1 _06013_ (.A(\tx_fifo.read_ptr[2] ),
    .Y(_00598_));
 sky130_fd_sc_hs__xnor2_1 _06014_ (.A(\tx_fifo.write_ptr[2] ),
    .B(_00598_),
    .Y(_00599_));
 sky130_fd_sc_hs__inv_1 _06015_ (.A(\tx_fifo.read_ptr[3] ),
    .Y(_00600_));
 sky130_fd_sc_hs__xnor2_1 _06016_ (.A(\tx_fifo.write_ptr[3] ),
    .B(_00600_),
    .Y(_00601_));
 sky130_fd_sc_hs__or2_1 _06017_ (.A(_00599_),
    .B(_00601_),
    .X(_00602_));
 sky130_fd_sc_hs__inv_2 _06018_ (.A(\tx_fifo.read_ptr[6] ),
    .Y(_00603_));
 sky130_fd_sc_hs__xnor2_1 _06019_ (.A(\tx_fifo.write_ptr[6] ),
    .B(_00603_),
    .Y(_00604_));
 sky130_fd_sc_hs__inv_1 _06020_ (.A(_00604_),
    .Y(_00605_));
 sky130_fd_sc_hs__xnor2_1 _06021_ (.A(\tx_fifo.write_ptr[7] ),
    .B(\tx_fifo.read_ptr[7] ),
    .Y(_00606_));
 sky130_fd_sc_hs__nand2_1 _06022_ (.A(_00605_),
    .B(_00606_),
    .Y(_00607_));
 sky130_fd_sc_hs__inv_2 _06023_ (.A(\tx_fifo.read_ptr[1] ),
    .Y(_00231_));
 sky130_fd_sc_hs__xnor2_1 _06024_ (.A(\tx_fifo.write_ptr[1] ),
    .B(_00231_),
    .Y(_00608_));
 sky130_fd_sc_hs__inv_2 _06025_ (.A(\tx_fifo.read_ptr[0] ),
    .Y(_00230_));
 sky130_fd_sc_hs__xnor2_1 _06026_ (.A(\tx_fifo.write_ptr[0] ),
    .B(_00230_),
    .Y(_00609_));
 sky130_fd_sc_hs__or2_1 _06027_ (.A(_00608_),
    .B(_00609_),
    .X(_00610_));
 sky130_fd_sc_hs__nor4_1 _06028_ (.A(_00597_),
    .B(_00602_),
    .C(_00607_),
    .D(_00610_),
    .Y(_00611_));
 sky130_fd_sc_hs__inv_1 _06029_ (.A(net3316),
    .Y(_00612_));
 sky130_fd_sc_hs__inv_2 _06030_ (.A(\u_window_buffer.current_state[2] ),
    .Y(_00613_));
 sky130_fd_sc_hs__nor2_1 _06031_ (.A(\u_window_buffer.move_counter[23] ),
    .B(\u_window_buffer.move_counter[22] ),
    .Y(_00614_));
 sky130_fd_sc_hs__inv_1 _06032_ (.A(_00614_),
    .Y(_00615_));
 sky130_fd_sc_hs__nor2_1 _06033_ (.A(\u_window_buffer.move_counter[21] ),
    .B(\u_window_buffer.move_counter[20] ),
    .Y(_00616_));
 sky130_fd_sc_hs__inv_1 _06034_ (.A(_00616_),
    .Y(_00617_));
 sky130_fd_sc_hs__nor2_1 _06035_ (.A(\u_window_buffer.move_counter[25] ),
    .B(\u_window_buffer.move_counter[26] ),
    .Y(_00618_));
 sky130_fd_sc_hs__inv_1 _06036_ (.A(\u_window_buffer.move_counter[24] ),
    .Y(_00619_));
 sky130_fd_sc_hs__inv_1 _06037_ (.A(\u_window_buffer.move_counter[27] ),
    .Y(_00620_));
 sky130_fd_sc_hs__nand3_1 _06038_ (.A(_00618_),
    .B(_00619_),
    .C(_00620_),
    .Y(_00621_));
 sky130_fd_sc_hs__nor3_1 _06039_ (.A(_00615_),
    .B(_00617_),
    .C(_00621_),
    .Y(_00622_));
 sky130_fd_sc_hs__nor2_1 _06040_ (.A(\u_window_buffer.move_counter[19] ),
    .B(\u_window_buffer.move_counter[18] ),
    .Y(_00623_));
 sky130_fd_sc_hs__inv_2 _06041_ (.A(_00623_),
    .Y(_00624_));
 sky130_fd_sc_hs__nor2_1 _06042_ (.A(\u_window_buffer.move_counter[17] ),
    .B(\u_window_buffer.move_counter[16] ),
    .Y(_00625_));
 sky130_fd_sc_hs__inv_1 _06043_ (.A(_00625_),
    .Y(_00626_));
 sky130_fd_sc_hs__nor2_1 _06044_ (.A(_00624_),
    .B(_00626_),
    .Y(_00627_));
 sky130_fd_sc_hs__nor2_1 _06045_ (.A(\u_window_buffer.move_counter[29] ),
    .B(\u_window_buffer.move_counter[30] ),
    .Y(_00628_));
 sky130_fd_sc_hs__nor2_1 _06046_ (.A(\u_window_buffer.move_counter[28] ),
    .B(\u_window_buffer.move_counter[31] ),
    .Y(_00629_));
 sky130_fd_sc_hs__nand4_1 _06047_ (.A(_00622_),
    .B(_00627_),
    .C(_00628_),
    .D(_00629_),
    .Y(_00630_));
 sky130_fd_sc_hs__nor2_1 _06048_ (.A(\u_window_buffer.move_counter[11] ),
    .B(\u_window_buffer.move_counter[10] ),
    .Y(_00631_));
 sky130_fd_sc_hs__inv_1 _06049_ (.A(_00631_),
    .Y(_00632_));
 sky130_fd_sc_hs__nor2_1 _06050_ (.A(\u_window_buffer.move_counter[9] ),
    .B(\u_window_buffer.move_counter[8] ),
    .Y(_00633_));
 sky130_fd_sc_hs__inv_2 _06051_ (.A(_00633_),
    .Y(_00634_));
 sky130_fd_sc_hs__nor2_1 _06052_ (.A(_00632_),
    .B(_00634_),
    .Y(_00635_));
 sky130_fd_sc_hs__nor2_1 _06053_ (.A(\u_window_buffer.move_counter[15] ),
    .B(\u_window_buffer.move_counter[14] ),
    .Y(_00636_));
 sky130_fd_sc_hs__nor2_1 _06054_ (.A(\u_window_buffer.move_counter[13] ),
    .B(\u_window_buffer.move_counter[12] ),
    .Y(_00637_));
 sky130_fd_sc_hs__nand3_1 _06055_ (.A(_00635_),
    .B(_00636_),
    .C(_00637_),
    .Y(_00638_));
 sky130_fd_sc_hs__inv_1 _06056_ (.A(_00223_),
    .Y(_00639_));
 sky130_fd_sc_hs__nor2_1 _06057_ (.A(\u_window_buffer.move_counter[3] ),
    .B(\u_window_buffer.move_counter[2] ),
    .Y(_00640_));
 sky130_fd_sc_hs__inv_1 _06058_ (.A(_00640_),
    .Y(_00641_));
 sky130_fd_sc_hs__nor2_1 _06059_ (.A(_00639_),
    .B(_00641_),
    .Y(_00642_));
 sky130_fd_sc_hs__inv_1 _06060_ (.A(_00642_),
    .Y(_00643_));
 sky130_fd_sc_hs__nor2_1 _06061_ (.A(\u_window_buffer.move_counter[5] ),
    .B(\u_window_buffer.move_counter[4] ),
    .Y(_00644_));
 sky130_fd_sc_hs__inv_1 _06062_ (.A(_00644_),
    .Y(_00645_));
 sky130_fd_sc_hs__nor2_1 _06063_ (.A(\u_window_buffer.move_counter[7] ),
    .B(\u_window_buffer.move_counter[6] ),
    .Y(_00646_));
 sky130_fd_sc_hs__inv_2 _06064_ (.A(_00646_),
    .Y(_00647_));
 sky130_fd_sc_hs__nor2_1 _06065_ (.A(_00645_),
    .B(_00647_),
    .Y(_00648_));
 sky130_fd_sc_hs__inv_1 _06066_ (.A(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hs__nor2_1 _06067_ (.A(_00643_),
    .B(_00649_),
    .Y(_00650_));
 sky130_fd_sc_hs__inv_1 _06068_ (.A(_00650_),
    .Y(_00651_));
 sky130_fd_sc_hs__nor2_1 _06069_ (.A(_00638_),
    .B(_00651_),
    .Y(_00652_));
 sky130_fd_sc_hs__inv_1 _06070_ (.A(_00652_),
    .Y(_00653_));
 sky130_fd_sc_hs__nor2_1 _06071_ (.A(_00630_),
    .B(_00653_),
    .Y(_00654_));
 sky130_fd_sc_hs__inv_1 _06072_ (.A(\u_window_buffer.current_state[4] ),
    .Y(_00655_));
 sky130_fd_sc_hs__o21ai_1 _06073_ (.A1(_00613_),
    .A2(_00654_),
    .B1(_00655_),
    .Y(_00656_));
 sky130_fd_sc_hs__clkinv_1 _06074_ (.A(_00656_),
    .Y(_00657_));
 sky130_fd_sc_hs__nor2_4 _06075_ (.A(\u_window_buffer.current_state[0] ),
    .B(\u_window_buffer.current_state[3] ),
    .Y(_00658_));
 sky130_fd_sc_hs__o21ai_1 _06076_ (.A1(_00612_),
    .A2(_00657_),
    .B1(_00658_),
    .Y(_00659_));
 sky130_fd_sc_hs__inv_2 _06077_ (.A(_00659_),
    .Y(_00660_));
 sky130_fd_sc_hs__nor2_1 _06078_ (.A(_05774_),
    .B(_00660_),
    .Y(_00021_));
 sky130_fd_sc_hs__or2_1 _06079_ (.A(_00006_),
    .B(_00021_),
    .X(_00024_));
 sky130_fd_sc_hs__nand2_1 _06080_ (.A(_00660_),
    .B(net3784),
    .Y(_00023_));
 sky130_fd_sc_hs__nor3_1 _06081_ (.A(net3782),
    .B(net3316),
    .C(_00657_),
    .Y(_00020_));
 sky130_fd_sc_hs__buf_1 place2187 (.A(_03453_),
    .X(net2187));
 sky130_fd_sc_hs__buf_1 place2186 (.A(_03467_),
    .X(net2186));
 sky130_fd_sc_hs__nand2_1 _06084_ (.A(_00654_),
    .B(\u_window_buffer.current_state[2] ),
    .Y(_00663_));
 sky130_fd_sc_hs__nor2_1 _06085_ (.A(start_move),
    .B(_00592_),
    .Y(_00664_));
 sky130_fd_sc_hs__inv_1 _06086_ (.A(_00664_),
    .Y(_00665_));
 sky130_fd_sc_hs__buf_1 place2185 (.A(_04537_),
    .X(net2185));
 sky130_fd_sc_hs__a21oi_1 _06088_ (.A1(_00663_),
    .A2(_00665_),
    .B1(net3782),
    .Y(_00019_));
 sky130_fd_sc_hs__a21oi_1 _06089_ (.A1(fft_done),
    .A2(\u_mel.state[0] ),
    .B1(mel_valid),
    .Y(_00667_));
 sky130_fd_sc_hs__nor2_1 _06090_ (.A(_00667_),
    .B(_05820_),
    .Y(_00017_));
 sky130_fd_sc_hs__a21oi_1 _06091_ (.A1(_00566_),
    .A2(\u_hamming_window.hamming_state[0] ),
    .B1(net3782),
    .Y(_00668_));
 sky130_fd_sc_hs__inv_2 _06092_ (.A(\u_hamming_window.hamming_state[3] ),
    .Y(_00669_));
 sky130_fd_sc_hs__nand2_1 _06093_ (.A(_00668_),
    .B(_00669_),
    .Y(_00012_));
 sky130_fd_sc_hs__inv_2 _06094_ (.A(net3744),
    .Y(_00150_));
 sky130_fd_sc_hs__inv_1 _06095_ (.A(_00148_),
    .Y(_00151_));
 sky130_fd_sc_hs__nand2_1 _06096_ (.A(_00114_),
    .B(net3538),
    .Y(_00670_));
 sky130_fd_sc_hs__nand2_1 _06097_ (.A(net3535),
    .B(net3533),
    .Y(_00671_));
 sky130_fd_sc_hs__or2_2 _06098_ (.A(_00670_),
    .B(_00671_),
    .X(_00672_));
 sky130_fd_sc_hs__nand2_1 _06099_ (.A(net3525),
    .B(net3523),
    .Y(_00673_));
 sky130_fd_sc_hs__inv_1 _06100_ (.A(_00125_),
    .Y(_00674_));
 sky130_fd_sc_hs__nand2_4 _06101_ (.A(_00673_),
    .B(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hs__and2_4 _06102_ (.A(net3530),
    .B(net3528),
    .X(_00676_));
 sky130_fd_sc_hs__nand2_1 _06103_ (.A(_00122_),
    .B(_00123_),
    .Y(_00677_));
 sky130_fd_sc_hs__inv_1 _06104_ (.A(net3532),
    .Y(_00678_));
 sky130_fd_sc_hs__nand2_1 _06105_ (.A(_00677_),
    .B(_00678_),
    .Y(_00679_));
 sky130_fd_sc_hs__a21oi_4 _06106_ (.A1(_00675_),
    .A2(_00676_),
    .B1(_00679_),
    .Y(_00680_));
 sky130_fd_sc_hs__a21oi_1 _06107_ (.A1(_00118_),
    .A2(_00119_),
    .B1(net3537),
    .Y(_00681_));
 sky130_fd_sc_hs__a21oi_1 _06108_ (.A1(_00114_),
    .A2(_00115_),
    .B1(_00113_),
    .Y(_00682_));
 sky130_fd_sc_hs__o21ai_4 _06109_ (.A1(net3496),
    .A2(net3493),
    .B1(net3491),
    .Y(_00683_));
 sky130_fd_sc_hs__o21bai_1 _06110_ (.A1(net3420),
    .A2(_00680_),
    .B1_N(_00683_),
    .Y(_00684_));
 sky130_fd_sc_hs__nand2_1 _06111_ (.A(_00098_),
    .B(net3555),
    .Y(_00685_));
 sky130_fd_sc_hs__nand2_1 _06112_ (.A(net3553),
    .B(net3551),
    .Y(_00686_));
 sky130_fd_sc_hs__nor2_1 _06113_ (.A(_00685_),
    .B(_00686_),
    .Y(_00687_));
 sky130_fd_sc_hs__inv_1 _06114_ (.A(_00687_),
    .Y(_00688_));
 sky130_fd_sc_hs__nand2_1 _06115_ (.A(net3548),
    .B(net3546),
    .Y(_00689_));
 sky130_fd_sc_hs__nand2_1 _06116_ (.A(_00110_),
    .B(net3541),
    .Y(_00690_));
 sky130_fd_sc_hs__nor2_1 _06117_ (.A(_00689_),
    .B(_00690_),
    .Y(_00691_));
 sky130_fd_sc_hs__inv_1 _06118_ (.A(_00691_),
    .Y(_00692_));
 sky130_fd_sc_hs__nor2_2 _06119_ (.A(_00688_),
    .B(_00692_),
    .Y(_00693_));
 sky130_fd_sc_hs__a21oi_1 _06120_ (.A1(_00110_),
    .A2(net3543),
    .B1(net3545),
    .Y(_00694_));
 sky130_fd_sc_hs__a21oi_1 _06121_ (.A1(_00106_),
    .A2(net3547),
    .B1(net3550),
    .Y(_00695_));
 sky130_fd_sc_hs__o21ai_2 _06122_ (.A1(net3487),
    .A2(net3486),
    .B1(net3484),
    .Y(_00696_));
 sky130_fd_sc_hs__nand2_1 _06123_ (.A(_00696_),
    .B(net3416),
    .Y(_00697_));
 sky130_fd_sc_hs__a21o_1 _06124_ (.A1(_00098_),
    .A2(net3556),
    .B1(_00097_),
    .X(_00698_));
 sky130_fd_sc_hs__a21oi_1 _06125_ (.A1(_00102_),
    .A2(net3552),
    .B1(net3554),
    .Y(_00699_));
 sky130_fd_sc_hs__nor2_1 _06126_ (.A(net3490),
    .B(net3482),
    .Y(_00700_));
 sky130_fd_sc_hs__nor2_1 _06127_ (.A(_00698_),
    .B(_00700_),
    .Y(_00701_));
 sky130_fd_sc_hs__nand2_1 _06128_ (.A(_00697_),
    .B(_00701_),
    .Y(_00702_));
 sky130_fd_sc_hs__a21oi_2 _06129_ (.A1(_00684_),
    .A2(_00693_),
    .B1(_00702_),
    .Y(_00703_));
 sky130_fd_sc_hs__nand2_1 _06130_ (.A(_00142_),
    .B(_00143_),
    .Y(_00704_));
 sky130_fd_sc_hs__inv_1 _06131_ (.A(_00141_),
    .Y(_00705_));
 sky130_fd_sc_hs__nand2_1 _06132_ (.A(_00704_),
    .B(_00705_),
    .Y(_00706_));
 sky130_fd_sc_hs__bufbuf_8 place2184 (.A(_04559_),
    .X(net2184));
 sky130_fd_sc_hs__buf_1 place2183 (.A(_04565_),
    .X(net2183));
 sky130_fd_sc_hs__and2_1 _06135_ (.A(_00138_),
    .B(_00140_),
    .X(_00709_));
 sky130_fd_sc_hs__nand2_1 _06136_ (.A(_00706_),
    .B(_00709_),
    .Y(_00710_));
 sky130_fd_sc_hs__a21oi_1 _06137_ (.A1(_00138_),
    .A2(_00139_),
    .B1(_00137_),
    .Y(_00711_));
 sky130_fd_sc_hs__nand2_1 _06138_ (.A(_00710_),
    .B(_00711_),
    .Y(_00712_));
 sky130_fd_sc_hs__nand2_2 _06139_ (.A(_00132_),
    .B(_00130_),
    .Y(_00713_));
 sky130_fd_sc_hs__nand2_2 _06140_ (.A(_00134_),
    .B(net3789),
    .Y(_00714_));
 sky130_fd_sc_hs__nor2_2 _06141_ (.A(_00713_),
    .B(_00714_),
    .Y(_00715_));
 sky130_fd_sc_hs__nand2_1 _06142_ (.A(_00712_),
    .B(_00715_),
    .Y(_00716_));
 sky130_fd_sc_hs__nand2_1 _06143_ (.A(_00134_),
    .B(_00135_),
    .Y(_00717_));
 sky130_fd_sc_hs__inv_1 _06144_ (.A(net3514),
    .Y(_00718_));
 sky130_fd_sc_hs__nand2_1 _06145_ (.A(_00717_),
    .B(_00718_),
    .Y(_00719_));
 sky130_fd_sc_hs__and2_1 _06146_ (.A(_00130_),
    .B(_00132_),
    .X(_00720_));
 sky130_fd_sc_hs__nand2_1 _06147_ (.A(_00130_),
    .B(_00131_),
    .Y(_00721_));
 sky130_fd_sc_hs__inv_1 _06148_ (.A(net3519),
    .Y(_00722_));
 sky130_fd_sc_hs__nand2_1 _06149_ (.A(_00721_),
    .B(_00722_),
    .Y(_00723_));
 sky130_fd_sc_hs__a21oi_2 _06150_ (.A1(_00719_),
    .A2(_00720_),
    .B1(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hs__nand2_2 _06151_ (.A(_00138_),
    .B(_00140_),
    .Y(_00725_));
 sky130_fd_sc_hs__buf_4 place2181 (.A(_05445_),
    .X(net2181));
 sky130_fd_sc_hs__nand2_2 _06153_ (.A(_00142_),
    .B(_00144_),
    .Y(_00727_));
 sky130_fd_sc_hs__nor2_4 _06154_ (.A(_00727_),
    .B(_00725_),
    .Y(_00728_));
 sky130_fd_sc_hs__nand2_2 _06155_ (.A(_00146_),
    .B(_00147_),
    .Y(_00729_));
 sky130_fd_sc_hs__inv_1 _06156_ (.A(_00145_),
    .Y(_00730_));
 sky130_fd_sc_hs__nand2_2 _06157_ (.A(_00730_),
    .B(_00729_),
    .Y(_00731_));
 sky130_fd_sc_hs__nand3_1 _06158_ (.A(net4875),
    .B(_00715_),
    .C(net3408),
    .Y(_00732_));
 sky130_fd_sc_hs__nand3_1 _06159_ (.A(_00716_),
    .B(_00724_),
    .C(_00732_),
    .Y(_00733_));
 sky130_fd_sc_hs__buf_1 place2182 (.A(net2181),
    .X(net2182));
 sky130_fd_sc_hs__and2_4 _06161_ (.A(net3527),
    .B(net3521),
    .X(_00735_));
 sky130_fd_sc_hs__nand2_2 _06162_ (.A(_00676_),
    .B(_00735_),
    .Y(_00736_));
 sky130_fd_sc_hs__nor2_4 _06163_ (.A(_00736_),
    .B(_00672_),
    .Y(_00737_));
 sky130_fd_sc_hs__nand3_2 _06164_ (.A(net3237),
    .B(_00693_),
    .C(net3356),
    .Y(_00738_));
 sky130_fd_sc_hs__nand2_2 _06165_ (.A(_00703_),
    .B(_00738_),
    .Y(_00739_));
 sky130_fd_sc_hs__inv_1 _06166_ (.A(_00090_),
    .Y(_00740_));
 sky130_fd_sc_hs__clkinv_1 _06167_ (.A(_00092_),
    .Y(_00741_));
 sky130_fd_sc_hs__inv_2 _06168_ (.A(_00094_),
    .Y(_00742_));
 sky130_fd_sc_hs__inv_1 _06169_ (.A(_00096_),
    .Y(_00743_));
 sky130_fd_sc_hs__nor2_1 _06170_ (.A(_00742_),
    .B(_00743_),
    .Y(_00744_));
 sky130_fd_sc_hs__inv_2 _06171_ (.A(_00744_),
    .Y(_00745_));
 sky130_fd_sc_hs__nor3_1 _06172_ (.A(_00740_),
    .B(_00741_),
    .C(net3355),
    .Y(_00746_));
 sky130_fd_sc_hs__nand2_1 _06173_ (.A(_00739_),
    .B(_00746_),
    .Y(_00747_));
 sky130_fd_sc_hs__nand2_1 _06174_ (.A(net3561),
    .B(net3560),
    .Y(_00748_));
 sky130_fd_sc_hs__inv_2 _06175_ (.A(_00093_),
    .Y(_00749_));
 sky130_fd_sc_hs__nand2_1 _06176_ (.A(_00748_),
    .B(_00749_),
    .Y(_00750_));
 sky130_fd_sc_hs__a21oi_1 _06177_ (.A1(net3404),
    .A2(net3563),
    .B1(_00091_),
    .Y(_00751_));
 sky130_fd_sc_hs__nor2_1 _06178_ (.A(net3476),
    .B(_00751_),
    .Y(_00752_));
 sky130_fd_sc_hs__nor2_1 _06179_ (.A(_00089_),
    .B(_00752_),
    .Y(_00753_));
 sky130_fd_sc_hs__nand2_1 _06180_ (.A(_00747_),
    .B(_00753_),
    .Y(_00754_));
 sky130_fd_sc_hs__xnor2_1 _06181_ (.A(\u_window_buffer.internal_read_ptr[31] ),
    .B(\u_window_buffer.read_ptr[31] ),
    .Y(_00755_));
 sky130_fd_sc_hs__inv_1 _06182_ (.A(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hs__nand2_1 _06183_ (.A(_00754_),
    .B(_00756_),
    .Y(_00757_));
 sky130_fd_sc_hs__nand3_1 _06184_ (.A(_00747_),
    .B(_00753_),
    .C(_00755_),
    .Y(_00758_));
 sky130_fd_sc_hs__and2_4 _06185_ (.A(_00758_),
    .B(_00757_),
    .X(_00759_));
 sky130_fd_sc_hs__bufbuf_8 place2180 (.A(_01686_),
    .X(net2180));
 sky130_fd_sc_hs__buf_1 place2179 (.A(_01704_),
    .X(net2179));
 sky130_fd_sc_hs__inv_4 _06188_ (.A(net2965),
    .Y(_00762_));
 sky130_fd_sc_hs__buf_1 place2178 (.A(_01714_),
    .X(net2178));
 sky130_fd_sc_hs__clkbuf_2 place2177 (.A(_03440_),
    .X(net2177));
 sky130_fd_sc_hs__nor2_1 _06191_ (.A(net3504),
    .B(net2966),
    .Y(_00765_));
 sky130_fd_sc_hs__inv_1 _06192_ (.A(_00765_),
    .Y(_00766_));
 sky130_fd_sc_hs__o21ai_1 _06193_ (.A1(_00153_),
    .A2(net2945),
    .B1(_00766_),
    .Y(_00154_));
 sky130_fd_sc_hs__bufbuf_8 place2176 (.A(_04549_),
    .X(net2176));
 sky130_fd_sc_hs__nand2_1 _06195_ (.A(_00138_),
    .B(net3510),
    .Y(_00768_));
 sky130_fd_sc_hs__inv_1 _06196_ (.A(_00137_),
    .Y(_00769_));
 sky130_fd_sc_hs__nand2_1 _06197_ (.A(_00768_),
    .B(_00769_),
    .Y(_00770_));
 sky130_fd_sc_hs__and2_1 _06198_ (.A(_00134_),
    .B(_00136_),
    .X(_00771_));
 sky130_fd_sc_hs__nand2_1 _06199_ (.A(_00770_),
    .B(_00771_),
    .Y(_00772_));
 sky130_fd_sc_hs__a21oi_1 _06200_ (.A1(_00134_),
    .A2(_00135_),
    .B1(net3515),
    .Y(_00773_));
 sky130_fd_sc_hs__nand2_1 _06201_ (.A(_00772_),
    .B(_00773_),
    .Y(_00774_));
 sky130_fd_sc_hs__inv_1 _06202_ (.A(_00774_),
    .Y(_00775_));
 sky130_fd_sc_hs__and2_1 _06203_ (.A(_00142_),
    .B(_00144_),
    .X(_00776_));
 sky130_fd_sc_hs__nand2_2 _06204_ (.A(_00731_),
    .B(_00776_),
    .Y(_00777_));
 sky130_fd_sc_hs__a21oi_1 _06205_ (.A1(_00142_),
    .A2(_00143_),
    .B1(_00141_),
    .Y(_00778_));
 sky130_fd_sc_hs__nand2_2 _06206_ (.A(_00777_),
    .B(_00778_),
    .Y(_00779_));
 sky130_fd_sc_hs__nor2_4 _06207_ (.A(_00714_),
    .B(_00725_),
    .Y(_00780_));
 sky130_fd_sc_hs__nand2_2 _06208_ (.A(_00779_),
    .B(_00780_),
    .Y(_00781_));
 sky130_fd_sc_hs__nand2_2 _06209_ (.A(_00781_),
    .B(_00775_),
    .Y(_00782_));
 sky130_fd_sc_hs__nand2_1 _06210_ (.A(net3521),
    .B(net3527),
    .Y(_00783_));
 sky130_fd_sc_hs__and2_1 _06211_ (.A(net3535),
    .B(net3533),
    .X(_00784_));
 sky130_fd_sc_hs__nand2_2 _06212_ (.A(_00676_),
    .B(_00784_),
    .Y(_00785_));
 sky130_fd_sc_hs__nor3_2 _06213_ (.A(_00783_),
    .B(net3480),
    .C(_00785_),
    .Y(_00786_));
 sky130_fd_sc_hs__nand2_1 _06214_ (.A(_00782_),
    .B(net3353),
    .Y(_00787_));
 sky130_fd_sc_hs__nand2_1 _06215_ (.A(net3419),
    .B(net3470),
    .Y(_00788_));
 sky130_fd_sc_hs__nand2_1 _06216_ (.A(_00788_),
    .B(net3494),
    .Y(_00789_));
 sky130_fd_sc_hs__a21oi_4 _06217_ (.A1(net3411),
    .A2(_00735_),
    .B1(_00675_),
    .Y(_00790_));
 sky130_fd_sc_hs__nor2_1 _06218_ (.A(net3403),
    .B(_00790_),
    .Y(_00791_));
 sky130_fd_sc_hs__nor2_1 _06219_ (.A(_00789_),
    .B(_00791_),
    .Y(_00792_));
 sky130_fd_sc_hs__nand2_1 _06220_ (.A(_00787_),
    .B(_00792_),
    .Y(_00793_));
 sky130_fd_sc_hs__nand2_1 _06221_ (.A(_00793_),
    .B(net3539),
    .Y(_00794_));
 sky130_fd_sc_hs__inv_1 _06222_ (.A(net3539),
    .Y(_00795_));
 sky130_fd_sc_hs__nand3_1 _06223_ (.A(net3193),
    .B(_00792_),
    .C(_00795_),
    .Y(_00796_));
 sky130_fd_sc_hs__nand2_2 _06224_ (.A(_00794_),
    .B(_00796_),
    .Y(_00797_));
 sky130_fd_sc_hs__nand2_1 _06225_ (.A(_00132_),
    .B(_00133_),
    .Y(_00798_));
 sky130_fd_sc_hs__inv_1 _06226_ (.A(_00131_),
    .Y(_00799_));
 sky130_fd_sc_hs__nand2_1 _06227_ (.A(_00798_),
    .B(_00799_),
    .Y(_00800_));
 sky130_fd_sc_hs__and2_1 _06228_ (.A(_00128_),
    .B(_00130_),
    .X(_00801_));
 sky130_fd_sc_hs__nand2_1 _06229_ (.A(_00800_),
    .B(_00801_),
    .Y(_00802_));
 sky130_fd_sc_hs__a21oi_1 _06230_ (.A1(_00128_),
    .A2(net3520),
    .B1(net3524),
    .Y(_00803_));
 sky130_fd_sc_hs__nand2_1 _06231_ (.A(_00802_),
    .B(_00803_),
    .Y(_00804_));
 sky130_fd_sc_hs__nand2_2 _06232_ (.A(_00120_),
    .B(_00122_),
    .Y(_00805_));
 sky130_fd_sc_hs__nand2_1 _06233_ (.A(_00124_),
    .B(_00126_),
    .Y(_00806_));
 sky130_fd_sc_hs__nor2_1 _06234_ (.A(net3469),
    .B(net3468),
    .Y(_00807_));
 sky130_fd_sc_hs__nand2_1 _06235_ (.A(_00124_),
    .B(_00125_),
    .Y(_00808_));
 sky130_fd_sc_hs__nand2b_1 _06236_ (.A_N(_00123_),
    .B(_00808_),
    .Y(_00809_));
 sky130_fd_sc_hs__inv_1 _06237_ (.A(_00805_),
    .Y(_00810_));
 sky130_fd_sc_hs__nand2_1 _06238_ (.A(_00809_),
    .B(net3401),
    .Y(_00811_));
 sky130_fd_sc_hs__nand2_1 _06239_ (.A(_00120_),
    .B(_00121_),
    .Y(_00812_));
 sky130_fd_sc_hs__inv_2 _06240_ (.A(_00119_),
    .Y(_00813_));
 sky130_fd_sc_hs__nand2_1 _06241_ (.A(_00812_),
    .B(_00813_),
    .Y(_00814_));
 sky130_fd_sc_hs__inv_1 _06242_ (.A(net3400),
    .Y(_00815_));
 sky130_fd_sc_hs__nand2_1 _06243_ (.A(_00811_),
    .B(_00815_),
    .Y(_00816_));
 sky130_fd_sc_hs__a21oi_1 _06244_ (.A1(_00804_),
    .A2(_00807_),
    .B1(_00816_),
    .Y(_00817_));
 sky130_fd_sc_hs__nand2_1 _06245_ (.A(_00140_),
    .B(_00141_),
    .Y(_00818_));
 sky130_fd_sc_hs__inv_1 _06246_ (.A(_00139_),
    .Y(_00819_));
 sky130_fd_sc_hs__nand2_1 _06247_ (.A(_00818_),
    .B(_00819_),
    .Y(_00820_));
 sky130_fd_sc_hs__and2_1 _06248_ (.A(_00138_),
    .B(_00136_),
    .X(_00821_));
 sky130_fd_sc_hs__nand2_1 _06249_ (.A(_00136_),
    .B(_00137_),
    .Y(_00822_));
 sky130_fd_sc_hs__inv_1 _06250_ (.A(_00135_),
    .Y(_00823_));
 sky130_fd_sc_hs__nand2_2 _06251_ (.A(_00822_),
    .B(_00823_),
    .Y(_00824_));
 sky130_fd_sc_hs__a21oi_4 _06252_ (.A1(_00820_),
    .A2(_00821_),
    .B1(net3399),
    .Y(_00825_));
 sky130_fd_sc_hs__a21oi_4 _06253_ (.A1(_00144_),
    .A2(_00145_),
    .B1(_00143_),
    .Y(_00826_));
 sky130_fd_sc_hs__nand3_2 _06254_ (.A(_00146_),
    .B(_00149_),
    .C(_00144_),
    .Y(_00827_));
 sky130_fd_sc_hs__nand2_2 _06255_ (.A(_00826_),
    .B(_00827_),
    .Y(_00828_));
 sky130_fd_sc_hs__nand2_1 _06256_ (.A(_00140_),
    .B(_00142_),
    .Y(_00829_));
 sky130_fd_sc_hs__nand2_1 _06257_ (.A(_00138_),
    .B(_00136_),
    .Y(_00830_));
 sky130_fd_sc_hs__nor2_2 _06258_ (.A(_00829_),
    .B(_00830_),
    .Y(_00831_));
 sky130_fd_sc_hs__nand2_2 _06259_ (.A(net4926),
    .B(_00831_),
    .Y(_00832_));
 sky130_fd_sc_hs__nand2_2 _06260_ (.A(_00832_),
    .B(_00825_),
    .Y(_00833_));
 sky130_fd_sc_hs__nand2_2 _06261_ (.A(_00128_),
    .B(_00130_),
    .Y(_00834_));
 sky130_fd_sc_hs__nand2_2 _06262_ (.A(_00134_),
    .B(_00132_),
    .Y(_00835_));
 sky130_fd_sc_hs__and2_1 _06263_ (.A(_00124_),
    .B(_00126_),
    .X(_00836_));
 sky130_fd_sc_hs__nand2_2 _06264_ (.A(_00810_),
    .B(_00836_),
    .Y(_00837_));
 sky130_fd_sc_hs__nor3_4 _06265_ (.A(net3465),
    .B(net3463),
    .C(net3350),
    .Y(_00838_));
 sky130_fd_sc_hs__nand2_2 _06266_ (.A(_00833_),
    .B(_00838_),
    .Y(_00839_));
 sky130_fd_sc_hs__nand2_1 _06267_ (.A(_00817_),
    .B(_00839_),
    .Y(_00840_));
 sky130_fd_sc_hs__inv_1 _06268_ (.A(net3536),
    .Y(_00841_));
 sky130_fd_sc_hs__nand2_2 _06269_ (.A(_00840_),
    .B(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hs__nand3_2 _06270_ (.A(net3271),
    .B(_00839_),
    .C(net3536),
    .Y(_00843_));
 sky130_fd_sc_hs__and2_1 _06271_ (.A(_00842_),
    .B(_00843_),
    .X(_00844_));
 sky130_fd_sc_hs__nand2_2 _06272_ (.A(_00797_),
    .B(_00844_),
    .Y(_00845_));
 sky130_fd_sc_hs__nand2_1 _06273_ (.A(_00144_),
    .B(net3506),
    .Y(_00846_));
 sky130_fd_sc_hs__inv_1 _06274_ (.A(_00143_),
    .Y(_00847_));
 sky130_fd_sc_hs__nand2_1 _06275_ (.A(_00846_),
    .B(_00847_),
    .Y(_00848_));
 sky130_fd_sc_hs__and2_2 _06276_ (.A(_00140_),
    .B(_00142_),
    .X(_00849_));
 sky130_fd_sc_hs__nand2_1 _06277_ (.A(_00848_),
    .B(_00849_),
    .Y(_00850_));
 sky130_fd_sc_hs__a21oi_2 _06278_ (.A1(_00140_),
    .A2(_00141_),
    .B1(_00139_),
    .Y(_00851_));
 sky130_fd_sc_hs__nand2_1 _06279_ (.A(_00850_),
    .B(_00851_),
    .Y(_00852_));
 sky130_fd_sc_hs__nor2_4 _06280_ (.A(_00835_),
    .B(_00830_),
    .Y(_00853_));
 sky130_fd_sc_hs__nand2_1 _06281_ (.A(_00852_),
    .B(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hs__inv_2 _06282_ (.A(_00835_),
    .Y(_00855_));
 sky130_fd_sc_hs__a21oi_4 _06283_ (.A1(_00824_),
    .A2(_00855_),
    .B1(_00800_),
    .Y(_00856_));
 sky130_fd_sc_hs__nand2_1 _06284_ (.A(net3505),
    .B(_00144_),
    .Y(_00857_));
 sky130_fd_sc_hs__nor2_1 _06285_ (.A(_00857_),
    .B(_00829_),
    .Y(_00858_));
 sky130_fd_sc_hs__nand3_2 _06286_ (.A(_00858_),
    .B(_00853_),
    .C(net3503),
    .Y(_00859_));
 sky130_fd_sc_hs__nand3_2 _06287_ (.A(_00859_),
    .B(_00856_),
    .C(_00854_),
    .Y(_00860_));
 sky130_fd_sc_hs__nand2_1 _06288_ (.A(_00116_),
    .B(_00118_),
    .Y(_00861_));
 sky130_fd_sc_hs__nor2_2 _06289_ (.A(_00805_),
    .B(_00861_),
    .Y(_00862_));
 sky130_fd_sc_hs__inv_1 _06290_ (.A(_00862_),
    .Y(_00863_));
 sky130_fd_sc_hs__nor3_4 _06291_ (.A(net3465),
    .B(net3468),
    .C(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hs__nand2_1 _06292_ (.A(net3235),
    .B(net3310),
    .Y(_00865_));
 sky130_fd_sc_hs__nand2_1 _06293_ (.A(_00128_),
    .B(_00129_),
    .Y(_00866_));
 sky130_fd_sc_hs__inv_1 _06294_ (.A(_00127_),
    .Y(_00867_));
 sky130_fd_sc_hs__nand2_1 _06295_ (.A(_00866_),
    .B(_00867_),
    .Y(_00868_));
 sky130_fd_sc_hs__nand2_1 _06296_ (.A(_00868_),
    .B(_00836_),
    .Y(_00869_));
 sky130_fd_sc_hs__a21oi_1 _06297_ (.A1(_00124_),
    .A2(_00125_),
    .B1(_00123_),
    .Y(_00870_));
 sky130_fd_sc_hs__nand2_1 _06298_ (.A(_00869_),
    .B(_00870_),
    .Y(_00871_));
 sky130_fd_sc_hs__nand2_1 _06299_ (.A(_00871_),
    .B(_00862_),
    .Y(_00872_));
 sky130_fd_sc_hs__clkinv_1 _06300_ (.A(_00861_),
    .Y(_00873_));
 sky130_fd_sc_hs__nand2_1 _06301_ (.A(_00873_),
    .B(_00814_),
    .Y(_00874_));
 sky130_fd_sc_hs__a21oi_1 _06302_ (.A1(_00116_),
    .A2(_00117_),
    .B1(_00115_),
    .Y(_00875_));
 sky130_fd_sc_hs__and2_1 _06303_ (.A(_00874_),
    .B(_00875_),
    .X(_00876_));
 sky130_fd_sc_hs__nand2_2 _06304_ (.A(_00872_),
    .B(_00876_),
    .Y(_00877_));
 sky130_fd_sc_hs__inv_1 _06305_ (.A(net3234),
    .Y(_00878_));
 sky130_fd_sc_hs__nand2_1 _06306_ (.A(_00865_),
    .B(_00878_),
    .Y(_00879_));
 sky130_fd_sc_hs__nand2_1 _06307_ (.A(_00879_),
    .B(net3540),
    .Y(_00880_));
 sky130_fd_sc_hs__inv_1 _06308_ (.A(net3540),
    .Y(_00881_));
 sky130_fd_sc_hs__nand3_1 _06309_ (.A(net3192),
    .B(_00881_),
    .C(net3191),
    .Y(_00882_));
 sky130_fd_sc_hs__nand2_2 _06310_ (.A(_00880_),
    .B(_00882_),
    .Y(_00883_));
 sky130_fd_sc_hs__nand2_1 _06311_ (.A(net3274),
    .B(net3359),
    .Y(_00884_));
 sky130_fd_sc_hs__nand2_1 _06312_ (.A(_00884_),
    .B(net3357),
    .Y(_00885_));
 sky130_fd_sc_hs__nor2_1 _06313_ (.A(_00672_),
    .B(_00680_),
    .Y(_00886_));
 sky130_fd_sc_hs__nor2_2 _06314_ (.A(net3417),
    .B(_00886_),
    .Y(_00887_));
 sky130_fd_sc_hs__inv_1 _06315_ (.A(net3542),
    .Y(_00888_));
 sky130_fd_sc_hs__nand4_1 _06316_ (.A(_00737_),
    .B(net3409),
    .C(net3410),
    .D(net3413),
    .Y(_00889_));
 sky130_fd_sc_hs__nand4_1 _06317_ (.A(net3190),
    .B(_00887_),
    .C(_00888_),
    .D(_00889_),
    .Y(_00890_));
 sky130_fd_sc_hs__nand3_1 _06318_ (.A(_00885_),
    .B(_00887_),
    .C(_00889_),
    .Y(_00891_));
 sky130_fd_sc_hs__nand2_1 _06319_ (.A(_00891_),
    .B(net3542),
    .Y(_00892_));
 sky130_fd_sc_hs__nand2_2 _06320_ (.A(_00892_),
    .B(_00890_),
    .Y(_00893_));
 sky130_fd_sc_hs__nand3b_2 _06321_ (.A_N(_00845_),
    .B(_00893_),
    .C(_00883_),
    .Y(_00894_));
 sky130_fd_sc_hs__nand2_2 _06322_ (.A(_00833_),
    .B(net3513),
    .Y(_00895_));
 sky130_fd_sc_hs__inv_1 _06323_ (.A(net3513),
    .Y(_00896_));
 sky130_fd_sc_hs__nand3_1 _06324_ (.A(_00825_),
    .B(net3352),
    .C(_00896_),
    .Y(_00897_));
 sky130_fd_sc_hs__and2_1 _06325_ (.A(_00895_),
    .B(_00897_),
    .X(_00898_));
 sky130_fd_sc_hs__inv_1 _06326_ (.A(net3516),
    .Y(_00899_));
 sky130_fd_sc_hs__nand2_1 _06327_ (.A(_00782_),
    .B(_00899_),
    .Y(_00900_));
 sky130_fd_sc_hs__nand3_1 _06328_ (.A(net3273),
    .B(net3272),
    .C(net3516),
    .Y(_00901_));
 sky130_fd_sc_hs__nand2_2 _06329_ (.A(_00901_),
    .B(_00900_),
    .Y(_00902_));
 sky130_fd_sc_hs__inv_1 _06330_ (.A(net3509),
    .Y(_00903_));
 sky130_fd_sc_hs__nand2_2 _06331_ (.A(_00779_),
    .B(_00903_),
    .Y(_00904_));
 sky130_fd_sc_hs__nand3_1 _06332_ (.A(net3354),
    .B(net3509),
    .C(net3471),
    .Y(_00905_));
 sky130_fd_sc_hs__nand2_2 _06333_ (.A(_00905_),
    .B(_00904_),
    .Y(_00906_));
 sky130_fd_sc_hs__nand2_1 _06334_ (.A(_00828_),
    .B(net3508),
    .Y(_00907_));
 sky130_fd_sc_hs__inv_1 _06335_ (.A(net3508),
    .Y(_00908_));
 sky130_fd_sc_hs__nand3_1 _06336_ (.A(net3467),
    .B(_00908_),
    .C(net3466),
    .Y(_00909_));
 sky130_fd_sc_hs__nand2_2 _06337_ (.A(_00907_),
    .B(_00909_),
    .Y(_00910_));
 sky130_fd_sc_hs__xnor2_2 _06338_ (.A(_00146_),
    .B(_00149_),
    .Y(_00911_));
 sky130_fd_sc_hs__nand2_1 _06339_ (.A(_00911_),
    .B(_00152_),
    .Y(_00912_));
 sky130_fd_sc_hs__inv_1 _06340_ (.A(net3507),
    .Y(_00913_));
 sky130_fd_sc_hs__nand2_1 _06341_ (.A(_00731_),
    .B(_00913_),
    .Y(_00914_));
 sky130_fd_sc_hs__nand3_1 _06342_ (.A(net4925),
    .B(net3477),
    .C(net3507),
    .Y(_00915_));
 sky130_fd_sc_hs__nand2_2 _06343_ (.A(_00914_),
    .B(_00915_),
    .Y(_00916_));
 sky130_fd_sc_hs__nor2_4 _06344_ (.A(_00916_),
    .B(_00912_),
    .Y(_00917_));
 sky130_fd_sc_hs__nand2_2 _06345_ (.A(_00910_),
    .B(_00917_),
    .Y(_00918_));
 sky130_fd_sc_hs__nor2_4 _06346_ (.A(_00918_),
    .B(_00906_),
    .Y(_00919_));
 sky130_fd_sc_hs__nand2_2 _06347_ (.A(_00828_),
    .B(net3462),
    .Y(_00920_));
 sky130_fd_sc_hs__nand2_1 _06348_ (.A(_00920_),
    .B(net3461),
    .Y(_00921_));
 sky130_fd_sc_hs__nand2_1 _06349_ (.A(_00921_),
    .B(net3511),
    .Y(_00922_));
 sky130_fd_sc_hs__inv_1 _06350_ (.A(net3511),
    .Y(_00923_));
 sky130_fd_sc_hs__nand3_1 _06351_ (.A(net3347),
    .B(_00923_),
    .C(net3461),
    .Y(_00924_));
 sky130_fd_sc_hs__nand2_2 _06352_ (.A(_00922_),
    .B(_00924_),
    .Y(_00925_));
 sky130_fd_sc_hs__nand2_2 _06353_ (.A(_00731_),
    .B(_00728_),
    .Y(_00926_));
 sky130_fd_sc_hs__nand3_2 _06354_ (.A(net3481),
    .B(_00710_),
    .C(_00926_),
    .Y(_00927_));
 sky130_fd_sc_hs__nand2_1 _06355_ (.A(_00927_),
    .B(net3512),
    .Y(_00928_));
 sky130_fd_sc_hs__inv_1 _06356_ (.A(net3512),
    .Y(_00929_));
 sky130_fd_sc_hs__nand4_1 _06357_ (.A(net3346),
    .B(net3360),
    .C(_00929_),
    .D(net3481),
    .Y(_00930_));
 sky130_fd_sc_hs__nand2_2 _06358_ (.A(_00930_),
    .B(_00928_),
    .Y(_00931_));
 sky130_fd_sc_hs__nand3_2 _06359_ (.A(_00931_),
    .B(_00925_),
    .C(_00919_),
    .Y(_00932_));
 sky130_fd_sc_hs__nor3_4 _06360_ (.A(_00932_),
    .B(_00902_),
    .C(_00898_),
    .Y(_00933_));
 sky130_fd_sc_hs__inv_1 _06361_ (.A(net3518),
    .Y(_00934_));
 sky130_fd_sc_hs__nand2_1 _06362_ (.A(_00860_),
    .B(_00934_),
    .Y(_00935_));
 sky130_fd_sc_hs__nand4_1 _06363_ (.A(_00854_),
    .B(net3349),
    .C(net3518),
    .D(_00859_),
    .Y(_00936_));
 sky130_fd_sc_hs__nand2_4 _06364_ (.A(_00935_),
    .B(_00936_),
    .Y(_00937_));
 sky130_fd_sc_hs__inv_1 _06365_ (.A(net3522),
    .Y(_00938_));
 sky130_fd_sc_hs__nand2_1 _06366_ (.A(net3237),
    .B(_00938_),
    .Y(_00939_));
 sky130_fd_sc_hs__nand4_1 _06367_ (.A(net3274),
    .B(net3359),
    .C(net3522),
    .D(net3358),
    .Y(_00940_));
 sky130_fd_sc_hs__nand2_2 _06368_ (.A(_00939_),
    .B(_00940_),
    .Y(_00941_));
 sky130_fd_sc_hs__nor2_4 _06369_ (.A(_00941_),
    .B(_00937_),
    .Y(_00942_));
 sky130_fd_sc_hs__nand2_1 _06370_ (.A(_00824_),
    .B(net3397),
    .Y(_00943_));
 sky130_fd_sc_hs__a21oi_1 _06371_ (.A1(_00132_),
    .A2(net3514),
    .B1(net3517),
    .Y(_00944_));
 sky130_fd_sc_hs__nand2_1 _06372_ (.A(_00943_),
    .B(_00944_),
    .Y(_00945_));
 sky130_fd_sc_hs__nor2_1 _06373_ (.A(_00834_),
    .B(_00806_),
    .Y(_00946_));
 sky130_fd_sc_hs__a21oi_2 _06374_ (.A1(_00945_),
    .A2(net3393),
    .B1(net3309),
    .Y(_00947_));
 sky130_fd_sc_hs__nand2_1 _06375_ (.A(net4905),
    .B(_00946_),
    .Y(_00948_));
 sky130_fd_sc_hs__clkinv_1 _06376_ (.A(_00948_),
    .Y(_00949_));
 sky130_fd_sc_hs__nand2_1 _06377_ (.A(net3306),
    .B(_00949_),
    .Y(_00950_));
 sky130_fd_sc_hs__nand2_1 _06378_ (.A(_00947_),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hs__inv_1 _06379_ (.A(net3531),
    .Y(_00952_));
 sky130_fd_sc_hs__nand2_1 _06380_ (.A(_00951_),
    .B(_00952_),
    .Y(_00953_));
 sky130_fd_sc_hs__nand3_1 _06381_ (.A(_00947_),
    .B(_00950_),
    .C(net3531),
    .Y(_00954_));
 sky130_fd_sc_hs__nand2_2 _06382_ (.A(_00953_),
    .B(_00954_),
    .Y(_00955_));
 sky130_fd_sc_hs__inv_1 _06383_ (.A(net3411),
    .Y(_00956_));
 sky130_fd_sc_hs__nand2_1 _06384_ (.A(net3412),
    .B(_00720_),
    .Y(_00957_));
 sky130_fd_sc_hs__nand2_1 _06385_ (.A(_00956_),
    .B(_00957_),
    .Y(_00958_));
 sky130_fd_sc_hs__inv_2 _06386_ (.A(net3406),
    .Y(_00959_));
 sky130_fd_sc_hs__a21o_1 _06387_ (.A1(_00675_),
    .A2(_00676_),
    .B1(_00679_),
    .X(_00960_));
 sky130_fd_sc_hs__a21oi_1 _06388_ (.A1(_00958_),
    .A2(_00959_),
    .B1(_00960_),
    .Y(_00961_));
 sky130_fd_sc_hs__nor3_4 _06389_ (.A(net3480),
    .B(net3478),
    .C(net3406),
    .Y(_00962_));
 sky130_fd_sc_hs__nand2_1 _06390_ (.A(_00927_),
    .B(_00962_),
    .Y(_00963_));
 sky130_fd_sc_hs__nand2_1 _06391_ (.A(_00961_),
    .B(_00963_),
    .Y(_00964_));
 sky130_fd_sc_hs__inv_1 _06392_ (.A(net3534),
    .Y(_00965_));
 sky130_fd_sc_hs__nand2_1 _06393_ (.A(_00964_),
    .B(_00965_),
    .Y(_00966_));
 sky130_fd_sc_hs__nand3_2 _06394_ (.A(net3269),
    .B(net3534),
    .C(_00963_),
    .Y(_00967_));
 sky130_fd_sc_hs__nand2_2 _06395_ (.A(_00966_),
    .B(_00967_),
    .Y(_00968_));
 sky130_fd_sc_hs__nor2_2 _06396_ (.A(_00955_),
    .B(_00968_),
    .Y(_00969_));
 sky130_fd_sc_hs__inv_1 _06397_ (.A(_00824_),
    .Y(_00970_));
 sky130_fd_sc_hs__nand2_1 _06398_ (.A(_00820_),
    .B(_00821_),
    .Y(_00971_));
 sky130_fd_sc_hs__nand2_1 _06399_ (.A(_00970_),
    .B(_00971_),
    .Y(_00972_));
 sky130_fd_sc_hs__nor2_2 _06400_ (.A(net3464),
    .B(_00835_),
    .Y(_00973_));
 sky130_fd_sc_hs__nand2_1 _06401_ (.A(_00972_),
    .B(_00973_),
    .Y(_00974_));
 sky130_fd_sc_hs__and2_2 _06402_ (.A(_00831_),
    .B(_00973_),
    .X(_00975_));
 sky130_fd_sc_hs__nand2_1 _06403_ (.A(_00975_),
    .B(net3791),
    .Y(_00976_));
 sky130_fd_sc_hs__a21oi_4 _06404_ (.A1(_00800_),
    .A2(_00801_),
    .B1(net3394),
    .Y(_00977_));
 sky130_fd_sc_hs__nand3_2 _06405_ (.A(_00974_),
    .B(_00976_),
    .C(net4877),
    .Y(_00978_));
 sky130_fd_sc_hs__inv_1 _06406_ (.A(net3526),
    .Y(_00979_));
 sky130_fd_sc_hs__nand2_1 _06407_ (.A(_00978_),
    .B(_00979_),
    .Y(_00980_));
 sky130_fd_sc_hs__nand4_1 _06408_ (.A(_00974_),
    .B(_00976_),
    .C(net3526),
    .D(net3343),
    .Y(_00981_));
 sky130_fd_sc_hs__nand2_1 _06409_ (.A(_00980_),
    .B(_00981_),
    .Y(_00982_));
 sky130_fd_sc_hs__nor2_2 _06410_ (.A(net3479),
    .B(_00783_),
    .Y(_00983_));
 sky130_fd_sc_hs__nand2_1 _06411_ (.A(_00774_),
    .B(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hs__and2_2 _06412_ (.A(_00983_),
    .B(_00780_),
    .X(_00985_));
 sky130_fd_sc_hs__nand2_2 _06413_ (.A(_00779_),
    .B(_00985_),
    .Y(_00986_));
 sky130_fd_sc_hs__nand3_2 _06414_ (.A(_00984_),
    .B(_00986_),
    .C(_00790_),
    .Y(_00987_));
 sky130_fd_sc_hs__nor2_2 _06415_ (.A(net3529),
    .B(_00987_),
    .Y(_00988_));
 sky130_fd_sc_hs__and2_2 _06416_ (.A(_00987_),
    .B(net3529),
    .X(_00989_));
 sky130_fd_sc_hs__nor2_1 _06417_ (.A(_00988_),
    .B(_00989_),
    .Y(_00990_));
 sky130_fd_sc_hs__nor2_2 _06418_ (.A(_00990_),
    .B(_00982_),
    .Y(_00991_));
 sky130_fd_sc_hs__nand4_2 _06419_ (.A(_00969_),
    .B(_00942_),
    .C(_00933_),
    .D(_00991_),
    .Y(_00992_));
 sky130_fd_sc_hs__nor2_4 _06420_ (.A(_00992_),
    .B(_00894_),
    .Y(_00993_));
 sky130_fd_sc_hs__nand2_1 _06421_ (.A(_00974_),
    .B(net3344),
    .Y(_00994_));
 sky130_fd_sc_hs__nand2_1 _06422_ (.A(_00112_),
    .B(_00114_),
    .Y(_00995_));
 sky130_fd_sc_hs__nor2_2 _06423_ (.A(_00861_),
    .B(_00995_),
    .Y(_00996_));
 sky130_fd_sc_hs__inv_2 _06424_ (.A(_00996_),
    .Y(_00997_));
 sky130_fd_sc_hs__nor2_2 _06425_ (.A(_00837_),
    .B(_00997_),
    .Y(_00998_));
 sky130_fd_sc_hs__nand2_1 _06426_ (.A(_00994_),
    .B(_00998_),
    .Y(_00999_));
 sky130_fd_sc_hs__a21oi_1 _06427_ (.A1(_00112_),
    .A2(_00113_),
    .B1(_00111_),
    .Y(_01000_));
 sky130_fd_sc_hs__o21ai_1 _06428_ (.A1(net3458),
    .A2(net3460),
    .B1(net3457),
    .Y(_01001_));
 sky130_fd_sc_hs__a21oi_4 _06429_ (.A1(net3314),
    .A2(net3392),
    .B1(_01001_),
    .Y(_01002_));
 sky130_fd_sc_hs__nand3_1 _06430_ (.A(_00998_),
    .B(net3398),
    .C(_00975_),
    .Y(_01003_));
 sky130_fd_sc_hs__nand3_1 _06431_ (.A(_00999_),
    .B(_01002_),
    .C(_01003_),
    .Y(_01004_));
 sky130_fd_sc_hs__nand2_1 _06432_ (.A(_01004_),
    .B(net3544),
    .Y(_01005_));
 sky130_fd_sc_hs__inv_1 _06433_ (.A(net3544),
    .Y(_01006_));
 sky130_fd_sc_hs__nand4_1 _06434_ (.A(_00999_),
    .B(_01002_),
    .C(_01003_),
    .D(_01006_),
    .Y(_01007_));
 sky130_fd_sc_hs__nand2_1 _06435_ (.A(_01005_),
    .B(_01007_),
    .Y(_01008_));
 sky130_fd_sc_hs__nand2_1 _06436_ (.A(net3268),
    .B(_00790_),
    .Y(_01009_));
 sky130_fd_sc_hs__or2_2 _06437_ (.A(_00690_),
    .B(net3495),
    .X(_01010_));
 sky130_fd_sc_hs__nor2_2 _06438_ (.A(_00785_),
    .B(_01010_),
    .Y(_01011_));
 sky130_fd_sc_hs__nand2_1 _06439_ (.A(_01009_),
    .B(_01011_),
    .Y(_01012_));
 sky130_fd_sc_hs__inv_2 _06440_ (.A(_01010_),
    .Y(_01013_));
 sky130_fd_sc_hs__o21ai_1 _06441_ (.A1(_00690_),
    .A2(net3492),
    .B1(net3486),
    .Y(_01014_));
 sky130_fd_sc_hs__a21oi_1 _06442_ (.A1(_00789_),
    .A2(_01013_),
    .B1(_01014_),
    .Y(_01015_));
 sky130_fd_sc_hs__nand3_1 _06443_ (.A(net3315),
    .B(_01011_),
    .C(net3342),
    .Y(_01016_));
 sky130_fd_sc_hs__nand3_1 _06444_ (.A(_01012_),
    .B(_01015_),
    .C(_01016_),
    .Y(_01017_));
 sky130_fd_sc_hs__nand2_1 _06445_ (.A(_01017_),
    .B(net3546),
    .Y(_01018_));
 sky130_fd_sc_hs__inv_1 _06446_ (.A(net3546),
    .Y(_01019_));
 sky130_fd_sc_hs__nand4_1 _06447_ (.A(_01012_),
    .B(_01015_),
    .C(_01016_),
    .D(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hs__nand2_1 _06448_ (.A(_01018_),
    .B(_01020_),
    .Y(_01021_));
 sky130_fd_sc_hs__nand2_1 _06449_ (.A(_01008_),
    .B(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hs__clkinv_1 _06450_ (.A(_01022_),
    .Y(_01023_));
 sky130_fd_sc_hs__o21ai_1 _06451_ (.A1(net3407),
    .A2(net3359),
    .B1(net3361),
    .Y(_01024_));
 sky130_fd_sc_hs__nor2_2 _06452_ (.A(net3420),
    .B(_00692_),
    .Y(_01025_));
 sky130_fd_sc_hs__nand2_1 _06453_ (.A(_01024_),
    .B(_01025_),
    .Y(_01026_));
 sky130_fd_sc_hs__a21oi_1 _06454_ (.A1(net3418),
    .A2(net3415),
    .B1(net3414),
    .Y(_01027_));
 sky130_fd_sc_hs__nand3_1 _06455_ (.A(net3305),
    .B(net3345),
    .C(_01025_),
    .Y(_01028_));
 sky130_fd_sc_hs__nand3_1 _06456_ (.A(_01026_),
    .B(_01027_),
    .C(_01028_),
    .Y(_01029_));
 sky130_fd_sc_hs__nand2_1 _06457_ (.A(_01029_),
    .B(net3551),
    .Y(_01030_));
 sky130_fd_sc_hs__inv_1 _06458_ (.A(net3551),
    .Y(_01031_));
 sky130_fd_sc_hs__nand4_1 _06459_ (.A(_01026_),
    .B(_01031_),
    .C(_01027_),
    .D(net3267),
    .Y(_01032_));
 sky130_fd_sc_hs__nand2_1 _06460_ (.A(_01030_),
    .B(_01032_),
    .Y(_01033_));
 sky130_fd_sc_hs__nand2_1 _06461_ (.A(_00945_),
    .B(net3393),
    .Y(_01034_));
 sky130_fd_sc_hs__a21oi_1 _06462_ (.A1(net3395),
    .A2(_00836_),
    .B1(net3402),
    .Y(_01035_));
 sky130_fd_sc_hs__nand2_1 _06463_ (.A(_01034_),
    .B(_01035_),
    .Y(_01036_));
 sky130_fd_sc_hs__nand2_1 _06464_ (.A(_00108_),
    .B(_00110_),
    .Y(_01037_));
 sky130_fd_sc_hs__nor2_2 _06465_ (.A(_01037_),
    .B(_00995_),
    .Y(_01038_));
 sky130_fd_sc_hs__nand2_1 _06466_ (.A(net3396),
    .B(_01038_),
    .Y(_01039_));
 sky130_fd_sc_hs__inv_1 _06467_ (.A(_01039_),
    .Y(_01040_));
 sky130_fd_sc_hs__nand2_1 _06468_ (.A(_01036_),
    .B(_01040_),
    .Y(_01041_));
 sky130_fd_sc_hs__nand2_1 _06469_ (.A(net3348),
    .B(net3460),
    .Y(_01042_));
 sky130_fd_sc_hs__a21oi_1 _06470_ (.A1(_00108_),
    .A2(_00109_),
    .B1(_00107_),
    .Y(_01043_));
 sky130_fd_sc_hs__o21ai_1 _06471_ (.A1(_01037_),
    .A2(_01000_),
    .B1(_01043_),
    .Y(_01044_));
 sky130_fd_sc_hs__a21oi_2 _06472_ (.A1(_01042_),
    .A2(_01038_),
    .B1(net3391),
    .Y(_01045_));
 sky130_fd_sc_hs__nor2_1 _06473_ (.A(_00948_),
    .B(_01039_),
    .Y(_01046_));
 sky130_fd_sc_hs__nand2_1 _06474_ (.A(net3306),
    .B(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hs__nand3_1 _06475_ (.A(_01041_),
    .B(_01045_),
    .C(_01047_),
    .Y(_01048_));
 sky130_fd_sc_hs__nand2_1 _06476_ (.A(_01048_),
    .B(net3549),
    .Y(_01049_));
 sky130_fd_sc_hs__inv_1 _06477_ (.A(net3549),
    .Y(_01050_));
 sky130_fd_sc_hs__nand4_1 _06478_ (.A(net3184),
    .B(_01045_),
    .C(_01050_),
    .D(_01047_),
    .Y(_01051_));
 sky130_fd_sc_hs__nand2_2 _06479_ (.A(_01049_),
    .B(_01051_),
    .Y(_01052_));
 sky130_fd_sc_hs__and2_1 _06480_ (.A(_01033_),
    .B(_01052_),
    .X(_01053_));
 sky130_fd_sc_hs__and2_1 _06481_ (.A(_01023_),
    .B(_01053_),
    .X(_01054_));
 sky130_fd_sc_hs__nand2_1 _06482_ (.A(_00993_),
    .B(_01054_),
    .Y(_01055_));
 sky130_fd_sc_hs__nand2_2 _06483_ (.A(_01055_),
    .B(_00759_),
    .Y(_01056_));
 sky130_fd_sc_hs__nor3_2 _06484_ (.A(net3488),
    .B(net3487),
    .C(_01010_),
    .Y(_01057_));
 sky130_fd_sc_hs__o21ai_1 _06485_ (.A1(_00789_),
    .A2(_00791_),
    .B1(_01057_),
    .Y(_01058_));
 sky130_fd_sc_hs__nor2_1 _06486_ (.A(net3489),
    .B(net3487),
    .Y(_01059_));
 sky130_fd_sc_hs__o21ai_1 _06487_ (.A1(net3489),
    .A2(net3485),
    .B1(net3482),
    .Y(_01060_));
 sky130_fd_sc_hs__a21oi_1 _06488_ (.A1(_01014_),
    .A2(_01059_),
    .B1(_01060_),
    .Y(_01061_));
 sky130_fd_sc_hs__and2_1 _06489_ (.A(_01057_),
    .B(net3353),
    .X(_01062_));
 sky130_fd_sc_hs__nand2_1 _06490_ (.A(_01062_),
    .B(net3236),
    .Y(_01063_));
 sky130_fd_sc_hs__nand3_1 _06491_ (.A(_01058_),
    .B(_01061_),
    .C(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hs__nand2_1 _06492_ (.A(_01064_),
    .B(net3555),
    .Y(_01065_));
 sky130_fd_sc_hs__inv_1 _06493_ (.A(net3555),
    .Y(_01066_));
 sky130_fd_sc_hs__nand4_1 _06494_ (.A(_01058_),
    .B(_01063_),
    .C(_01061_),
    .D(_01066_),
    .Y(_01067_));
 sky130_fd_sc_hs__nand2_1 _06495_ (.A(_01065_),
    .B(_01067_),
    .Y(_01068_));
 sky130_fd_sc_hs__o21bai_1 _06496_ (.A1(net3351),
    .A2(net3344),
    .B1_N(net3313),
    .Y(_01069_));
 sky130_fd_sc_hs__nand2_1 _06497_ (.A(_00106_),
    .B(_00104_),
    .Y(_01070_));
 sky130_fd_sc_hs__nor2_2 _06498_ (.A(net3456),
    .B(_01070_),
    .Y(_01071_));
 sky130_fd_sc_hs__inv_2 _06499_ (.A(_01071_),
    .Y(_01072_));
 sky130_fd_sc_hs__nor2_1 _06500_ (.A(_01072_),
    .B(net3341),
    .Y(_01073_));
 sky130_fd_sc_hs__nand2_1 _06501_ (.A(_01069_),
    .B(net3302),
    .Y(_01074_));
 sky130_fd_sc_hs__a21oi_1 _06502_ (.A1(_00104_),
    .A2(_00105_),
    .B1(_00103_),
    .Y(_01075_));
 sky130_fd_sc_hs__o21ai_1 _06503_ (.A1(net3454),
    .A2(net3455),
    .B1(net3453),
    .Y(_01076_));
 sky130_fd_sc_hs__a21oi_1 _06504_ (.A1(_01001_),
    .A2(_01071_),
    .B1(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hs__nand3_1 _06505_ (.A(net3312),
    .B(net3311),
    .C(net3302),
    .Y(_01078_));
 sky130_fd_sc_hs__nand3_1 _06506_ (.A(_01074_),
    .B(_01077_),
    .C(_01078_),
    .Y(_01079_));
 sky130_fd_sc_hs__nand2_1 _06507_ (.A(_01079_),
    .B(net3553),
    .Y(_01080_));
 sky130_fd_sc_hs__nand2_1 _06508_ (.A(_00840_),
    .B(net3303),
    .Y(_01081_));
 sky130_fd_sc_hs__inv_1 _06509_ (.A(net3553),
    .Y(_01082_));
 sky130_fd_sc_hs__nand3_1 _06510_ (.A(_01081_),
    .B(_01082_),
    .C(_01077_),
    .Y(_01083_));
 sky130_fd_sc_hs__nand2_1 _06511_ (.A(_01080_),
    .B(_01083_),
    .Y(_01084_));
 sky130_fd_sc_hs__nand2_2 _06512_ (.A(_01068_),
    .B(_01084_),
    .Y(_01085_));
 sky130_fd_sc_hs__nand2_1 _06513_ (.A(_00759_),
    .B(net2997),
    .Y(_01086_));
 sky130_fd_sc_hs__nand2_1 _06514_ (.A(_01056_),
    .B(_01086_),
    .Y(_01087_));
 sky130_fd_sc_hs__nand2_1 _06515_ (.A(_00100_),
    .B(_00102_),
    .Y(_01088_));
 sky130_fd_sc_hs__nor2_1 _06516_ (.A(_01088_),
    .B(_01070_),
    .Y(_01089_));
 sky130_fd_sc_hs__and2_1 _06517_ (.A(_01038_),
    .B(_01089_),
    .X(_01090_));
 sky130_fd_sc_hs__nand2_1 _06518_ (.A(_01044_),
    .B(_01089_),
    .Y(_01091_));
 sky130_fd_sc_hs__a21oi_1 _06519_ (.A1(_00100_),
    .A2(_00101_),
    .B1(_00099_),
    .Y(_01092_));
 sky130_fd_sc_hs__o21a_1 _06520_ (.A1(_01088_),
    .A2(_01075_),
    .B1(_01092_),
    .X(_01093_));
 sky130_fd_sc_hs__nand2_1 _06521_ (.A(_01091_),
    .B(_01093_),
    .Y(_01094_));
 sky130_fd_sc_hs__a21oi_1 _06522_ (.A1(_00877_),
    .A2(_01090_),
    .B1(_01094_),
    .Y(_01095_));
 sky130_fd_sc_hs__nand3_2 _06523_ (.A(_00860_),
    .B(net3310),
    .C(net3339),
    .Y(_01096_));
 sky130_fd_sc_hs__nand2_2 _06524_ (.A(net3182),
    .B(_01096_),
    .Y(_01097_));
 sky130_fd_sc_hs__nand2_1 _06525_ (.A(_01097_),
    .B(net3557),
    .Y(_01098_));
 sky130_fd_sc_hs__inv_1 _06526_ (.A(net3557),
    .Y(_01099_));
 sky130_fd_sc_hs__nand3_1 _06527_ (.A(net3183),
    .B(net3181),
    .C(_01099_),
    .Y(_01100_));
 sky130_fd_sc_hs__nand2_1 _06528_ (.A(_01098_),
    .B(_01100_),
    .Y(_01101_));
 sky130_fd_sc_hs__nand2_1 _06529_ (.A(_01087_),
    .B(net3039),
    .Y(_01102_));
 sky130_fd_sc_hs__and2_2 _06530_ (.A(_01098_),
    .B(_01100_),
    .X(_01103_));
 sky130_fd_sc_hs__nand3_1 _06531_ (.A(_01056_),
    .B(net3038),
    .C(_01086_),
    .Y(_01104_));
 sky130_fd_sc_hs__nand2_2 _06532_ (.A(_01104_),
    .B(_01102_),
    .Y(_01105_));
 sky130_fd_sc_hs__nand2_1 _06533_ (.A(_00739_),
    .B(net3473),
    .Y(_01106_));
 sky130_fd_sc_hs__nand3_1 _06534_ (.A(_00703_),
    .B(net3559),
    .C(_00738_),
    .Y(_01107_));
 sky130_fd_sc_hs__nand2_2 _06535_ (.A(_01106_),
    .B(_01107_),
    .Y(_01108_));
 sky130_fd_sc_hs__o31ai_2 _06536_ (.A1(_01103_),
    .A2(_01108_),
    .A3(_01085_),
    .B1(_00759_),
    .Y(_01109_));
 sky130_fd_sc_hs__nand2_1 _06537_ (.A(_01056_),
    .B(_01109_),
    .Y(_01110_));
 sky130_fd_sc_hs__nand2_1 _06538_ (.A(net3314),
    .B(net3392),
    .Y(_01111_));
 sky130_fd_sc_hs__o21a_1 _06539_ (.A1(net3458),
    .A2(net3460),
    .B1(net3457),
    .X(_01112_));
 sky130_fd_sc_hs__nand2_1 _06540_ (.A(_01111_),
    .B(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hs__nand2_1 _06541_ (.A(_00096_),
    .B(_00098_),
    .Y(_01114_));
 sky130_fd_sc_hs__nor3_4 _06542_ (.A(net3452),
    .B(_01114_),
    .C(_01072_),
    .Y(_01115_));
 sky130_fd_sc_hs__nor2_1 _06543_ (.A(net3452),
    .B(_01114_),
    .Y(_01116_));
 sky130_fd_sc_hs__nand2_1 _06544_ (.A(_01076_),
    .B(_01116_),
    .Y(_01117_));
 sky130_fd_sc_hs__a21oi_1 _06545_ (.A1(_00096_),
    .A2(net3558),
    .B1(_00095_),
    .Y(_01118_));
 sky130_fd_sc_hs__o21a_1 _06546_ (.A1(net3450),
    .A2(net3451),
    .B1(_01118_),
    .X(_01119_));
 sky130_fd_sc_hs__nand2_1 _06547_ (.A(_01117_),
    .B(_01119_),
    .Y(_01120_));
 sky130_fd_sc_hs__a21oi_4 _06548_ (.A1(_01113_),
    .A2(_01115_),
    .B1(_01120_),
    .Y(_01121_));
 sky130_fd_sc_hs__nand3_1 _06549_ (.A(_00978_),
    .B(net3304),
    .C(_01115_),
    .Y(_01122_));
 sky130_fd_sc_hs__nand2_1 _06550_ (.A(_01121_),
    .B(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hs__nand2_1 _06551_ (.A(_01123_),
    .B(net3474),
    .Y(_01124_));
 sky130_fd_sc_hs__nand3_1 _06552_ (.A(_01121_),
    .B(_01122_),
    .C(net3561),
    .Y(_01125_));
 sky130_fd_sc_hs__nand2_1 _06553_ (.A(_01124_),
    .B(_01125_),
    .Y(_01126_));
 sky130_fd_sc_hs__inv_1 _06554_ (.A(net3035),
    .Y(_01127_));
 sky130_fd_sc_hs__nand2_2 _06555_ (.A(_01110_),
    .B(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hs__nand2_1 _06556_ (.A(_01052_),
    .B(_01021_),
    .Y(_01129_));
 sky130_fd_sc_hs__nand2_2 _06557_ (.A(_01008_),
    .B(_00893_),
    .Y(_01130_));
 sky130_fd_sc_hs__nor2_4 _06558_ (.A(_01130_),
    .B(_01129_),
    .Y(_01131_));
 sky130_fd_sc_hs__or2_1 _06559_ (.A(net3186),
    .B(net3185),
    .X(_01132_));
 sky130_fd_sc_hs__and2_1 _06560_ (.A(net3188),
    .B(net3228),
    .X(_01133_));
 sky130_fd_sc_hs__nand2_1 _06561_ (.A(_01132_),
    .B(_01133_),
    .Y(_01134_));
 sky130_fd_sc_hs__nor2_2 _06562_ (.A(_00941_),
    .B(_00982_),
    .Y(_01135_));
 sky130_fd_sc_hs__nor2_1 _06563_ (.A(_00902_),
    .B(_00937_),
    .Y(_01136_));
 sky130_fd_sc_hs__nand2_1 _06564_ (.A(_00895_),
    .B(_00897_),
    .Y(_01137_));
 sky130_fd_sc_hs__nand2_1 _06565_ (.A(_01137_),
    .B(net4870),
    .Y(_01138_));
 sky130_fd_sc_hs__nor2_1 _06566_ (.A(net3744),
    .B(_00148_),
    .Y(_01139_));
 sky130_fd_sc_hs__nand2_1 _06567_ (.A(_00911_),
    .B(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hs__nor2_1 _06568_ (.A(_01140_),
    .B(_00916_),
    .Y(_01141_));
 sky130_fd_sc_hs__nand2_1 _06569_ (.A(_00910_),
    .B(_01141_),
    .Y(_01142_));
 sky130_fd_sc_hs__nor2_2 _06570_ (.A(_00906_),
    .B(_01142_),
    .Y(_01143_));
 sky130_fd_sc_hs__nand2_1 _06571_ (.A(_01143_),
    .B(_00925_),
    .Y(_01144_));
 sky130_fd_sc_hs__nor2_4 _06572_ (.A(_01144_),
    .B(_01138_),
    .Y(_01145_));
 sky130_fd_sc_hs__nand3_1 _06573_ (.A(_01135_),
    .B(_01136_),
    .C(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hs__nor2_2 _06574_ (.A(_01134_),
    .B(_01146_),
    .Y(_01147_));
 sky130_fd_sc_hs__and2_1 _06575_ (.A(net3187),
    .B(net3227),
    .X(_01148_));
 sky130_fd_sc_hs__nand2_1 _06576_ (.A(_00883_),
    .B(_01148_),
    .Y(_01149_));
 sky130_fd_sc_hs__nor2_1 _06577_ (.A(net2999),
    .B(_01149_),
    .Y(_01150_));
 sky130_fd_sc_hs__nand3_2 _06578_ (.A(_01131_),
    .B(_01147_),
    .C(_01150_),
    .Y(_01151_));
 sky130_fd_sc_hs__nand2_1 _06579_ (.A(_01151_),
    .B(_00759_),
    .Y(_01152_));
 sky130_fd_sc_hs__nand2_2 _06580_ (.A(_01084_),
    .B(_01033_),
    .Y(_01153_));
 sky130_fd_sc_hs__nand2_2 _06581_ (.A(_01101_),
    .B(_01068_),
    .Y(_01154_));
 sky130_fd_sc_hs__or2_1 _06582_ (.A(_01153_),
    .B(_01154_),
    .X(_01155_));
 sky130_fd_sc_hs__nand2_1 _06583_ (.A(_00759_),
    .B(_01155_),
    .Y(_01156_));
 sky130_fd_sc_hs__nand3_1 _06584_ (.A(_01152_),
    .B(net3037),
    .C(_01156_),
    .Y(_01157_));
 sky130_fd_sc_hs__nand2_1 _06585_ (.A(_00842_),
    .B(_00843_),
    .Y(_01158_));
 sky130_fd_sc_hs__nor2_1 _06586_ (.A(_01158_),
    .B(net3139),
    .Y(_01159_));
 sky130_fd_sc_hs__nand3_2 _06587_ (.A(_01159_),
    .B(_00883_),
    .C(net3046),
    .Y(_01160_));
 sky130_fd_sc_hs__and2_2 _06588_ (.A(_01136_),
    .B(_01145_),
    .X(_01161_));
 sky130_fd_sc_hs__nor2_1 _06589_ (.A(_00955_),
    .B(_00990_),
    .Y(_01162_));
 sky130_fd_sc_hs__nand3_2 _06590_ (.A(_01161_),
    .B(_01162_),
    .C(net3092),
    .Y(_01163_));
 sky130_fd_sc_hs__nor2_4 _06591_ (.A(_01160_),
    .B(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hs__nor2_4 _06592_ (.A(_01153_),
    .B(_01154_),
    .Y(_01165_));
 sky130_fd_sc_hs__nand3_1 _06593_ (.A(_01164_),
    .B(net2962),
    .C(_01165_),
    .Y(_01166_));
 sky130_fd_sc_hs__inv_1 _06594_ (.A(net3037),
    .Y(_01167_));
 sky130_fd_sc_hs__nand3_1 _06595_ (.A(_01166_),
    .B(_00759_),
    .C(_01167_),
    .Y(_01168_));
 sky130_fd_sc_hs__and2_2 _06596_ (.A(_01157_),
    .B(_01168_),
    .X(_01169_));
 sky130_fd_sc_hs__nand3_2 _06597_ (.A(_01056_),
    .B(net3035),
    .C(_01109_),
    .Y(_01170_));
 sky130_fd_sc_hs__nand3_2 _06598_ (.A(_01128_),
    .B(_01169_),
    .C(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hs__nor2_2 _06599_ (.A(_01126_),
    .B(net3036),
    .Y(_01172_));
 sky130_fd_sc_hs__nand4_2 _06600_ (.A(_01165_),
    .B(_01164_),
    .C(net2962),
    .D(_01172_),
    .Y(_01173_));
 sky130_fd_sc_hs__nand2_1 _06601_ (.A(_01173_),
    .B(_00759_),
    .Y(_01174_));
 sky130_fd_sc_hs__nand2_1 _06602_ (.A(_00789_),
    .B(_01013_),
    .Y(_01175_));
 sky130_fd_sc_hs__nand2b_1 _06603_ (.A_N(_01014_),
    .B(_01175_),
    .Y(_01176_));
 sky130_fd_sc_hs__nor3_2 _06604_ (.A(net3487),
    .B(_00745_),
    .C(_00688_),
    .Y(_01177_));
 sky130_fd_sc_hs__nor2_1 _06605_ (.A(net3490),
    .B(_00745_),
    .Y(_01178_));
 sky130_fd_sc_hs__nand2_1 _06606_ (.A(_01178_),
    .B(_01060_),
    .Y(_01179_));
 sky130_fd_sc_hs__a21oi_1 _06607_ (.A1(net3483),
    .A2(net3405),
    .B1(_00750_),
    .Y(_01180_));
 sky130_fd_sc_hs__nand2_1 _06608_ (.A(_01179_),
    .B(_01180_),
    .Y(_01181_));
 sky130_fd_sc_hs__a21oi_1 _06609_ (.A1(_01176_),
    .A2(_01177_),
    .B1(_01181_),
    .Y(_01182_));
 sky130_fd_sc_hs__nand3_2 _06610_ (.A(net3226),
    .B(net3340),
    .C(_01177_),
    .Y(_01183_));
 sky130_fd_sc_hs__nand2_1 _06611_ (.A(_01182_),
    .B(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hs__nand2_1 _06612_ (.A(_01184_),
    .B(net3475),
    .Y(_01185_));
 sky130_fd_sc_hs__nand3_1 _06613_ (.A(_01182_),
    .B(_01183_),
    .C(net3562),
    .Y(_01186_));
 sky130_fd_sc_hs__nand2_1 _06614_ (.A(_01185_),
    .B(_01186_),
    .Y(_01187_));
 sky130_fd_sc_hs__inv_1 _06615_ (.A(net3031),
    .Y(_01188_));
 sky130_fd_sc_hs__nand2_1 _06616_ (.A(_01174_),
    .B(net2993),
    .Y(_01189_));
 sky130_fd_sc_hs__nand3_1 _06617_ (.A(_01173_),
    .B(_00759_),
    .C(net3031),
    .Y(_01190_));
 sky130_fd_sc_hs__nand2_2 _06618_ (.A(_01189_),
    .B(_01190_),
    .Y(_01191_));
 sky130_fd_sc_hs__and2_2 _06619_ (.A(_01080_),
    .B(_01083_),
    .X(_01192_));
 sky130_fd_sc_hs__and2_2 _06620_ (.A(_01065_),
    .B(_01067_),
    .X(_01193_));
 sky130_fd_sc_hs__nor2_1 _06621_ (.A(_01192_),
    .B(_01193_),
    .Y(_01194_));
 sky130_fd_sc_hs__nand2_1 _06622_ (.A(_01194_),
    .B(_01053_),
    .Y(_01195_));
 sky130_fd_sc_hs__nor2_1 _06623_ (.A(_01103_),
    .B(_01108_),
    .Y(_01196_));
 sky130_fd_sc_hs__nor2_1 _06624_ (.A(_01126_),
    .B(_01187_),
    .Y(_01197_));
 sky130_fd_sc_hs__nand2_1 _06625_ (.A(_01196_),
    .B(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hs__nor2_2 _06626_ (.A(_01195_),
    .B(_01198_),
    .Y(_01199_));
 sky130_fd_sc_hs__nand3_2 _06627_ (.A(_01199_),
    .B(net2943),
    .C(net2963),
    .Y(_01200_));
 sky130_fd_sc_hs__nand2_1 _06628_ (.A(_01200_),
    .B(net2967),
    .Y(_01201_));
 sky130_fd_sc_hs__nor3_1 _06629_ (.A(_00741_),
    .B(net3474),
    .C(net3449),
    .Y(_01202_));
 sky130_fd_sc_hs__nand2_1 _06630_ (.A(net3136),
    .B(_01202_),
    .Y(_01203_));
 sky130_fd_sc_hs__o21ai_1 _06631_ (.A1(net3474),
    .A2(net3448),
    .B1(net3472),
    .Y(_01204_));
 sky130_fd_sc_hs__a21oi_1 _06632_ (.A1(_01204_),
    .A2(_00092_),
    .B1(_00091_),
    .Y(_01205_));
 sky130_fd_sc_hs__nand2_1 _06633_ (.A(_01203_),
    .B(_01205_),
    .Y(_01206_));
 sky130_fd_sc_hs__xnor2_2 _06634_ (.A(net3564),
    .B(_01206_),
    .Y(_01207_));
 sky130_fd_sc_hs__nand2_1 _06635_ (.A(_01201_),
    .B(net2992),
    .Y(_01208_));
 sky130_fd_sc_hs__nand3b_1 _06636_ (.A_N(net2992),
    .B(_01200_),
    .C(net2967),
    .Y(_01209_));
 sky130_fd_sc_hs__nand2_2 _06637_ (.A(_01208_),
    .B(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hs__nor2_2 _06638_ (.A(_01191_),
    .B(_01210_),
    .Y(_01211_));
 sky130_fd_sc_hs__o21ai_4 _06639_ (.A1(_01105_),
    .A2(_01171_),
    .B1(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hs__nand3_1 _06640_ (.A(_00759_),
    .B(_01207_),
    .C(_01188_),
    .Y(_01213_));
 sky130_fd_sc_hs__nor2_1 _06641_ (.A(_01213_),
    .B(_01173_),
    .Y(_01214_));
 sky130_fd_sc_hs__nand2_1 _06642_ (.A(net2900),
    .B(_01214_),
    .Y(_01215_));
 sky130_fd_sc_hs__nand2_2 _06643_ (.A(_01212_),
    .B(_01215_),
    .Y(_01216_));
 sky130_fd_sc_hs__inv_2 _06644_ (.A(net2835),
    .Y(_01217_));
 sky130_fd_sc_hs__nand2_2 _06645_ (.A(_01216_),
    .B(_01217_),
    .Y(_01218_));
 sky130_fd_sc_hs__nand3_2 _06646_ (.A(_01212_),
    .B(net2835),
    .C(_01215_),
    .Y(_01219_));
 sky130_fd_sc_hs__nand3_1 _06647_ (.A(_01214_),
    .B(net2967),
    .C(net2930),
    .Y(_01220_));
 sky130_fd_sc_hs__and2_2 _06648_ (.A(_01220_),
    .B(net2868),
    .X(_01221_));
 sky130_fd_sc_hs__o21a_1 _06649_ (.A1(net3033),
    .A2(net2942),
    .B1(_00759_),
    .X(_01222_));
 sky130_fd_sc_hs__xnor2_1 _06650_ (.A(net3030),
    .B(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hs__nand4_4 _06651_ (.A(_01218_),
    .B(_01219_),
    .C(_01221_),
    .D(net2896),
    .Y(_01224_));
 sky130_fd_sc_hs__nand2_1 _06652_ (.A(_01128_),
    .B(net2867),
    .Y(_01225_));
 sky130_fd_sc_hs__nand2_2 _06653_ (.A(_01225_),
    .B(_01220_),
    .Y(_01226_));
 sky130_fd_sc_hs__nor3_4 _06654_ (.A(net2866),
    .B(_01216_),
    .C(_01226_),
    .Y(_01227_));
 sky130_fd_sc_hs__nand2_2 _06655_ (.A(_01227_),
    .B(_01224_),
    .Y(_01228_));
 sky130_fd_sc_hs__nand3b_1 _06656_ (.A_N(net2853),
    .B(_01212_),
    .C(net2899),
    .Y(_01229_));
 sky130_fd_sc_hs__nand2_2 _06657_ (.A(_01228_),
    .B(net2808),
    .Y(_01230_));
 sky130_fd_sc_hs__nand2_2 _06658_ (.A(_01230_),
    .B(net2898),
    .Y(_01231_));
 sky130_fd_sc_hs__inv_1 _06659_ (.A(net2897),
    .Y(_01232_));
 sky130_fd_sc_hs__nand3_2 _06660_ (.A(_01232_),
    .B(net4864),
    .C(net2808),
    .Y(_01233_));
 sky130_fd_sc_hs__xnor2_1 _06661_ (.A(net3091),
    .B(net2901),
    .Y(_01234_));
 sky130_fd_sc_hs__inv_1 _06662_ (.A(_01234_),
    .Y(_01235_));
 sky130_fd_sc_hs__nand2_2 _06663_ (.A(_01218_),
    .B(net2809),
    .Y(_01236_));
 sky130_fd_sc_hs__inv_1 _06664_ (.A(net2799),
    .Y(_01237_));
 sky130_fd_sc_hs__nand4_2 _06665_ (.A(_01231_),
    .B(_01233_),
    .C(_01235_),
    .D(_01237_),
    .Y(_01238_));
 sky130_fd_sc_hs__inv_1 _06666_ (.A(_01229_),
    .Y(_01239_));
 sky130_fd_sc_hs__o21ai_1 _06667_ (.A1(_01239_),
    .A2(_01227_),
    .B1(_01224_),
    .Y(_01240_));
 sky130_fd_sc_hs__nand2_1 _06668_ (.A(_01217_),
    .B(_01221_),
    .Y(_01241_));
 sky130_fd_sc_hs__xnor2_1 _06669_ (.A(_01226_),
    .B(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hs__and3_1 _06670_ (.A(_01212_),
    .B(_01226_),
    .C(_01215_),
    .X(_01243_));
 sky130_fd_sc_hs__a21oi_1 _06671_ (.A1(_01242_),
    .A2(_01216_),
    .B1(_01243_),
    .Y(_01244_));
 sky130_fd_sc_hs__inv_1 _06672_ (.A(net2798),
    .Y(_01245_));
 sky130_fd_sc_hs__nand2_1 _06673_ (.A(_01240_),
    .B(_01245_),
    .Y(_01246_));
 sky130_fd_sc_hs__o211ai_1 _06674_ (.A1(_01239_),
    .A2(_01227_),
    .B1(_01244_),
    .C1(_01224_),
    .Y(_01247_));
 sky130_fd_sc_hs__nand2_2 _06675_ (.A(_01246_),
    .B(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hs__inv_1 _06676_ (.A(_01221_),
    .Y(_01249_));
 sky130_fd_sc_hs__nor2_1 _06677_ (.A(net2869),
    .B(net2835),
    .Y(_01250_));
 sky130_fd_sc_hs__nor2_1 _06678_ (.A(_01217_),
    .B(_01249_),
    .Y(_01251_));
 sky130_fd_sc_hs__o21ai_1 _06679_ (.A1(_01250_),
    .A2(_01251_),
    .B1(net3792),
    .Y(_01252_));
 sky130_fd_sc_hs__o21ai_2 _06680_ (.A1(net2834),
    .A2(net4862),
    .B1(_01252_),
    .Y(_01253_));
 sky130_fd_sc_hs__o21ai_1 _06681_ (.A1(_01232_),
    .A2(_01236_),
    .B1(_01253_),
    .Y(_01254_));
 sky130_fd_sc_hs__nand4_1 _06682_ (.A(net2804),
    .B(net2810),
    .C(net2834),
    .D(net2896),
    .Y(_01255_));
 sky130_fd_sc_hs__nand2_1 _06683_ (.A(_01254_),
    .B(_01255_),
    .Y(_01256_));
 sky130_fd_sc_hs__nand2_1 _06684_ (.A(_01256_),
    .B(_01230_),
    .Y(_01257_));
 sky130_fd_sc_hs__nand3_1 _06685_ (.A(_01228_),
    .B(net2808),
    .C(_01253_),
    .Y(_01258_));
 sky130_fd_sc_hs__nand2_2 _06686_ (.A(_01257_),
    .B(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hs__nor2_2 _06687_ (.A(_01248_),
    .B(_01259_),
    .Y(_01260_));
 sky130_fd_sc_hs__nand2_2 _06688_ (.A(_01260_),
    .B(_01238_),
    .Y(_01261_));
 sky130_fd_sc_hs__o21ai_1 _06689_ (.A1(net2866),
    .A2(net2811),
    .B1(_01247_),
    .Y(_01262_));
 sky130_fd_sc_hs__nand2_2 _06690_ (.A(_01262_),
    .B(_01228_),
    .Y(_01263_));
 sky130_fd_sc_hs__nand2_2 _06691_ (.A(_01263_),
    .B(_01261_),
    .Y(_01264_));
 sky130_fd_sc_hs__nand2_1 _06692_ (.A(_01231_),
    .B(_01233_),
    .Y(_01265_));
 sky130_fd_sc_hs__xnor2_1 _06693_ (.A(net2898),
    .B(net2799),
    .Y(_01266_));
 sky130_fd_sc_hs__nand2_1 _06694_ (.A(net2781),
    .B(_01266_),
    .Y(_01267_));
 sky130_fd_sc_hs__o21ai_2 _06695_ (.A1(net2800),
    .A2(net2781),
    .B1(_01267_),
    .Y(_01268_));
 sky130_fd_sc_hs__o21ai_1 _06696_ (.A1(net2865),
    .A2(_01265_),
    .B1(_01268_),
    .Y(_01269_));
 sky130_fd_sc_hs__nand4_1 _06697_ (.A(net2774),
    .B(net2780),
    .C(net2852),
    .D(net2800),
    .Y(_01270_));
 sky130_fd_sc_hs__nand2_1 _06698_ (.A(_01269_),
    .B(_01270_),
    .Y(_01271_));
 sky130_fd_sc_hs__nand2_1 _06699_ (.A(_01264_),
    .B(_01271_),
    .Y(_01272_));
 sky130_fd_sc_hs__nand3_1 _06700_ (.A(_01261_),
    .B(_01268_),
    .C(_01263_),
    .Y(_01273_));
 sky130_fd_sc_hs__nand2_1 _06701_ (.A(_01272_),
    .B(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hs__nand3_1 _06702_ (.A(_01231_),
    .B(_01233_),
    .C(_01237_),
    .Y(_01275_));
 sky130_fd_sc_hs__nor2_1 _06703_ (.A(net2865),
    .B(_01275_),
    .Y(_01276_));
 sky130_fd_sc_hs__nand2_1 _06704_ (.A(_01276_),
    .B(net2763),
    .Y(_01277_));
 sky130_fd_sc_hs__inv_1 _06705_ (.A(_01259_),
    .Y(_01278_));
 sky130_fd_sc_hs__nand2_1 _06706_ (.A(net2765),
    .B(_01278_),
    .Y(_01279_));
 sky130_fd_sc_hs__nand2_1 _06707_ (.A(_01277_),
    .B(_01279_),
    .Y(_01280_));
 sky130_fd_sc_hs__nand2_2 _06708_ (.A(_01280_),
    .B(_01264_),
    .Y(_01281_));
 sky130_fd_sc_hs__nand3_1 _06709_ (.A(net2749),
    .B(net2772),
    .C(net2764),
    .Y(_01282_));
 sky130_fd_sc_hs__nand2_1 _06710_ (.A(_01281_),
    .B(_01282_),
    .Y(_01283_));
 sky130_fd_sc_hs__nor2_2 _06711_ (.A(_01283_),
    .B(_01274_),
    .Y(_01284_));
 sky130_fd_sc_hs__nand2_2 _06712_ (.A(net2852),
    .B(_01264_),
    .Y(_01285_));
 sky130_fd_sc_hs__xnor2_1 _06713_ (.A(net3137),
    .B(net2931),
    .Y(_01286_));
 sky130_fd_sc_hs__inv_1 _06714_ (.A(net2762),
    .Y(_01287_));
 sky130_fd_sc_hs__o211ai_2 _06715_ (.A1(_01248_),
    .A2(_01259_),
    .B1(net2865),
    .C1(_01263_),
    .Y(_01288_));
 sky130_fd_sc_hs__nand4_2 _06716_ (.A(_01285_),
    .B(net2894),
    .C(_01287_),
    .D(_01288_),
    .Y(_01289_));
 sky130_fd_sc_hs__nand2_2 _06717_ (.A(_01289_),
    .B(_01284_),
    .Y(_01290_));
 sky130_fd_sc_hs__nor2_1 _06718_ (.A(net2763),
    .B(_01276_),
    .Y(_01291_));
 sky130_fd_sc_hs__nand2_1 _06719_ (.A(_01264_),
    .B(_01291_),
    .Y(_01292_));
 sky130_fd_sc_hs__inv_1 _06720_ (.A(net2773),
    .Y(_01293_));
 sky130_fd_sc_hs__nand2_1 _06721_ (.A(_01292_),
    .B(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hs__nand3_1 _06722_ (.A(_01264_),
    .B(net2773),
    .C(_01291_),
    .Y(_01295_));
 sky130_fd_sc_hs__nand2_2 _06723_ (.A(_01294_),
    .B(_01295_),
    .Y(_01296_));
 sky130_fd_sc_hs__inv_2 _06724_ (.A(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hs__nand2_2 _06725_ (.A(_01297_),
    .B(_01290_),
    .Y(_01298_));
 sky130_fd_sc_hs__nand2_2 _06726_ (.A(_01298_),
    .B(net2895),
    .Y(_01299_));
 sky130_fd_sc_hs__inv_1 _06727_ (.A(net2894),
    .Y(_01300_));
 sky130_fd_sc_hs__nand3_2 _06728_ (.A(net2864),
    .B(_01290_),
    .C(_01297_),
    .Y(_01301_));
 sky130_fd_sc_hs__o31ai_1 _06729_ (.A1(net2998),
    .A2(net2964),
    .A3(net3043),
    .B1(net2965),
    .Y(_01302_));
 sky130_fd_sc_hs__xnor2_1 _06730_ (.A(net3040),
    .B(_01302_),
    .Y(_01303_));
 sky130_fd_sc_hs__nand2_2 _06731_ (.A(_01285_),
    .B(_01288_),
    .Y(_01304_));
 sky130_fd_sc_hs__inv_1 _06732_ (.A(net2725),
    .Y(_01305_));
 sky130_fd_sc_hs__nand4_2 _06733_ (.A(_01299_),
    .B(_01301_),
    .C(net2928),
    .D(_01305_),
    .Y(_01306_));
 sky130_fd_sc_hs__and2_1 _06734_ (.A(_01281_),
    .B(net2739),
    .X(_01307_));
 sky130_fd_sc_hs__inv_1 _06735_ (.A(net2727),
    .Y(_01308_));
 sky130_fd_sc_hs__o211ai_2 _06736_ (.A1(_01296_),
    .A2(_01307_),
    .B1(_01308_),
    .C1(net2726),
    .Y(_01309_));
 sky130_fd_sc_hs__a21o_1 _06737_ (.A1(net2726),
    .A2(_01296_),
    .B1(_01308_),
    .X(_01310_));
 sky130_fd_sc_hs__nand2_2 _06738_ (.A(_01309_),
    .B(_01310_),
    .Y(_01311_));
 sky130_fd_sc_hs__nand2_1 _06739_ (.A(_01285_),
    .B(net2762),
    .Y(_01312_));
 sky130_fd_sc_hs__nor2_1 _06740_ (.A(net2865),
    .B(net2762),
    .Y(_01313_));
 sky130_fd_sc_hs__nand2_1 _06741_ (.A(net3802),
    .B(_01313_),
    .Y(_01314_));
 sky130_fd_sc_hs__nand2_2 _06742_ (.A(_01312_),
    .B(_01314_),
    .Y(_01315_));
 sky130_fd_sc_hs__nor2_2 _06743_ (.A(_01300_),
    .B(_01304_),
    .Y(_01316_));
 sky130_fd_sc_hs__or2_1 _06744_ (.A(_01315_),
    .B(_01316_),
    .X(_01317_));
 sky130_fd_sc_hs__nand2_1 _06745_ (.A(_01316_),
    .B(_01315_),
    .Y(_01318_));
 sky130_fd_sc_hs__nand2_1 _06746_ (.A(_01317_),
    .B(_01318_),
    .Y(_01319_));
 sky130_fd_sc_hs__nand2_1 _06747_ (.A(_01319_),
    .B(_01298_),
    .Y(_01320_));
 sky130_fd_sc_hs__nand3b_1 _06748_ (.A_N(net2720),
    .B(_01290_),
    .C(net2708),
    .Y(_01321_));
 sky130_fd_sc_hs__nand2_2 _06749_ (.A(_01320_),
    .B(_01321_),
    .Y(_01322_));
 sky130_fd_sc_hs__nor2_2 _06750_ (.A(_01311_),
    .B(_01322_),
    .Y(_01323_));
 sky130_fd_sc_hs__nand2_2 _06751_ (.A(_01306_),
    .B(_01323_),
    .Y(_01324_));
 sky130_fd_sc_hs__inv_1 _06752_ (.A(net2709),
    .Y(_01325_));
 sky130_fd_sc_hs__a31oi_2 _06753_ (.A1(_01308_),
    .A2(net2726),
    .A3(_01296_),
    .B1(_01307_),
    .Y(_01326_));
 sky130_fd_sc_hs__or2_4 _06754_ (.A(_01326_),
    .B(_01325_),
    .X(_01327_));
 sky130_fd_sc_hs__nand2_2 _06755_ (.A(_01324_),
    .B(_01327_),
    .Y(_01328_));
 sky130_fd_sc_hs__nand2_2 _06756_ (.A(_01328_),
    .B(net2929),
    .Y(_01329_));
 sky130_fd_sc_hs__inv_1 _06757_ (.A(net2928),
    .Y(_01330_));
 sky130_fd_sc_hs__nand3_2 _06758_ (.A(net2690),
    .B(net2893),
    .C(_01324_),
    .Y(_01331_));
 sky130_fd_sc_hs__o31ai_1 _06759_ (.A1(net2996),
    .A2(net2995),
    .A3(net2994),
    .B1(net2965),
    .Y(_01332_));
 sky130_fd_sc_hs__xnor2_1 _06760_ (.A(net3041),
    .B(_01332_),
    .Y(_01333_));
 sky130_fd_sc_hs__and2_2 _06761_ (.A(_01299_),
    .B(_01301_),
    .X(_01334_));
 sky130_fd_sc_hs__nand4_2 _06762_ (.A(_01329_),
    .B(_01331_),
    .C(net2926),
    .D(net2678),
    .Y(_01335_));
 sky130_fd_sc_hs__and2_1 _06763_ (.A(_01309_),
    .B(_01310_),
    .X(_01336_));
 sky130_fd_sc_hs__nor2_1 _06764_ (.A(_01325_),
    .B(_01326_),
    .Y(_01337_));
 sky130_fd_sc_hs__clkinv_1 _06765_ (.A(_01322_),
    .Y(_01338_));
 sky130_fd_sc_hs__o211ai_2 _06766_ (.A1(_01336_),
    .A2(_01337_),
    .B1(_01338_),
    .C1(net3806),
    .Y(_01339_));
 sky130_fd_sc_hs__nand3_1 _06767_ (.A(_01299_),
    .B(_01301_),
    .C(_01305_),
    .Y(_01340_));
 sky130_fd_sc_hs__nor2_1 _06768_ (.A(_01330_),
    .B(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hs__o21ai_2 _06769_ (.A1(_01327_),
    .A2(_01341_),
    .B1(net2679),
    .Y(_01342_));
 sky130_fd_sc_hs__nand2_1 _06770_ (.A(_01339_),
    .B(_01342_),
    .Y(_01343_));
 sky130_fd_sc_hs__nand2_1 _06771_ (.A(_01334_),
    .B(net2929),
    .Y(_01344_));
 sky130_fd_sc_hs__nand2_1 _06772_ (.A(_01299_),
    .B(net2725),
    .Y(_01345_));
 sky130_fd_sc_hs__nand2_1 _06773_ (.A(net2699),
    .B(net2719),
    .Y(_01346_));
 sky130_fd_sc_hs__and2_2 _06774_ (.A(_01345_),
    .B(_01346_),
    .X(_01347_));
 sky130_fd_sc_hs__nand2_1 _06775_ (.A(_01344_),
    .B(_01347_),
    .Y(_01348_));
 sky130_fd_sc_hs__nand4_1 _06776_ (.A(net2691),
    .B(net2698),
    .C(net2928),
    .D(net2725),
    .Y(_01349_));
 sky130_fd_sc_hs__nand2_1 _06777_ (.A(_01348_),
    .B(_01349_),
    .Y(_01350_));
 sky130_fd_sc_hs__nand2_2 _06778_ (.A(_01328_),
    .B(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hs__nand3_1 _06779_ (.A(_01324_),
    .B(_01347_),
    .C(net2690),
    .Y(_01352_));
 sky130_fd_sc_hs__nand2_2 _06780_ (.A(_01351_),
    .B(_01352_),
    .Y(_01353_));
 sky130_fd_sc_hs__nor2_4 _06781_ (.A(_01343_),
    .B(_01353_),
    .Y(_01354_));
 sky130_fd_sc_hs__nand2_2 _06782_ (.A(_01335_),
    .B(_01354_),
    .Y(_01355_));
 sky130_fd_sc_hs__nand4_1 _06783_ (.A(net2681),
    .B(_01338_),
    .C(net2697),
    .D(net2689),
    .Y(_01356_));
 sky130_fd_sc_hs__o21ai_1 _06784_ (.A1(net2680),
    .A2(_01341_),
    .B1(net2696),
    .Y(_01357_));
 sky130_fd_sc_hs__nand2_1 _06785_ (.A(_01356_),
    .B(_01357_),
    .Y(_01358_));
 sky130_fd_sc_hs__inv_1 _06786_ (.A(_01358_),
    .Y(_01359_));
 sky130_fd_sc_hs__nand2_2 _06787_ (.A(_01355_),
    .B(_01359_),
    .Y(_01360_));
 sky130_fd_sc_hs__nand2_2 _06788_ (.A(_01360_),
    .B(net2927),
    .Y(_01361_));
 sky130_fd_sc_hs__o21ai_1 _06789_ (.A1(net2964),
    .A2(net3043),
    .B1(net2965),
    .Y(_01362_));
 sky130_fd_sc_hs__xnor2_1 _06790_ (.A(net3042),
    .B(_01362_),
    .Y(_01363_));
 sky130_fd_sc_hs__and2_2 _06791_ (.A(_01329_),
    .B(_01331_),
    .X(_01364_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _06792_ (.A(net2926),
    .Y(_01365_));
 sky130_fd_sc_hs__nand3b_4 _06793_ (.A_N(_01354_),
    .B(_01365_),
    .C(_01359_),
    .Y(_01366_));
 sky130_fd_sc_hs__nand4_2 _06794_ (.A(_01361_),
    .B(net2924),
    .C(net2632),
    .D(_01366_),
    .Y(_01367_));
 sky130_fd_sc_hs__o21ai_1 _06795_ (.A1(net2649),
    .A2(_01354_),
    .B1(net2636),
    .Y(_01368_));
 sky130_fd_sc_hs__nand2_1 _06796_ (.A(net2635),
    .B(_01368_),
    .Y(_01369_));
 sky130_fd_sc_hs__and2_1 _06797_ (.A(_01339_),
    .B(_01342_),
    .X(_01370_));
 sky130_fd_sc_hs__inv_1 _06798_ (.A(_01353_),
    .Y(_01371_));
 sky130_fd_sc_hs__o211ai_2 _06799_ (.A1(_01358_),
    .A2(_01370_),
    .B1(_01371_),
    .C1(_01335_),
    .Y(_01372_));
 sky130_fd_sc_hs__nand2_2 _06800_ (.A(_01369_),
    .B(_01372_),
    .Y(_01373_));
 sky130_fd_sc_hs__nand2_1 _06801_ (.A(net2691),
    .B(net2698),
    .Y(_01374_));
 sky130_fd_sc_hs__nand2_1 _06802_ (.A(net2643),
    .B(net2676),
    .Y(_01375_));
 sky130_fd_sc_hs__nor2_1 _06803_ (.A(net2893),
    .B(_01374_),
    .Y(_01376_));
 sky130_fd_sc_hs__nand2_1 _06804_ (.A(net2652),
    .B(_01376_),
    .Y(_01377_));
 sky130_fd_sc_hs__and2_2 _06805_ (.A(_01375_),
    .B(_01377_),
    .X(_01378_));
 sky130_fd_sc_hs__nand2_1 _06806_ (.A(_01364_),
    .B(net2927),
    .Y(_01379_));
 sky130_fd_sc_hs__nand2_1 _06807_ (.A(_01378_),
    .B(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hs__nand4_1 _06808_ (.A(net2643),
    .B(net2651),
    .C(net2927),
    .D(net2677),
    .Y(_01381_));
 sky130_fd_sc_hs__nand2_1 _06809_ (.A(_01380_),
    .B(_01381_),
    .Y(_01382_));
 sky130_fd_sc_hs__nand2_1 _06810_ (.A(_01360_),
    .B(_01382_),
    .Y(_01383_));
 sky130_fd_sc_hs__nand3_1 _06811_ (.A(_01355_),
    .B(_01359_),
    .C(_01378_),
    .Y(_01384_));
 sky130_fd_sc_hs__nand2_2 _06812_ (.A(_01383_),
    .B(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hs__nor2_4 _06813_ (.A(_01373_),
    .B(_01385_),
    .Y(_01386_));
 sky130_fd_sc_hs__nand2_2 _06814_ (.A(_01367_),
    .B(_01386_),
    .Y(_01387_));
 sky130_fd_sc_hs__nand2_1 _06815_ (.A(_01372_),
    .B(net2650),
    .Y(_01388_));
 sky130_fd_sc_hs__and2_2 _06816_ (.A(_01388_),
    .B(net3833),
    .X(_01389_));
 sky130_fd_sc_hs__clkinv_1 _06817_ (.A(_01389_),
    .Y(_01390_));
 sky130_fd_sc_hs__nand2_2 _06818_ (.A(_01390_),
    .B(_01387_),
    .Y(_01391_));
 sky130_fd_sc_hs__nand2_2 _06819_ (.A(_01391_),
    .B(net2925),
    .Y(_01392_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _06820_ (.A(net2923),
    .Y(_01393_));
 sky130_fd_sc_hs__nand3_2 _06821_ (.A(_01387_),
    .B(net2892),
    .C(net2596),
    .Y(_01394_));
 sky130_fd_sc_hs__nor2_1 _06822_ (.A(net2961),
    .B(_00762_),
    .Y(_01395_));
 sky130_fd_sc_hs__xnor2_1 _06823_ (.A(net3044),
    .B(_01395_),
    .Y(_01396_));
 sky130_fd_sc_hs__inv_1 _06824_ (.A(_01396_),
    .Y(_01397_));
 sky130_fd_sc_hs__and2_2 _06825_ (.A(net2607),
    .B(net2616),
    .X(_01398_));
 sky130_fd_sc_hs__nand4_4 _06826_ (.A(_01392_),
    .B(_01394_),
    .C(_01397_),
    .D(net2595),
    .Y(_01399_));
 sky130_fd_sc_hs__o21ai_1 _06827_ (.A1(net2604),
    .A2(_01386_),
    .B1(net2598),
    .Y(_01400_));
 sky130_fd_sc_hs__nand2_1 _06828_ (.A(_01400_),
    .B(net2597),
    .Y(_01401_));
 sky130_fd_sc_hs__and2_1 _06829_ (.A(net4872),
    .B(_01372_),
    .X(_01402_));
 sky130_fd_sc_hs__inv_1 _06830_ (.A(net2597),
    .Y(_01403_));
 sky130_fd_sc_hs__o211ai_1 _06831_ (.A1(_01402_),
    .A2(_01389_),
    .B1(net2599),
    .C1(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hs__nand2_1 _06832_ (.A(_01401_),
    .B(_01404_),
    .Y(_01405_));
 sky130_fd_sc_hs__nand2_1 _06833_ (.A(_01398_),
    .B(net2925),
    .Y(_01406_));
 sky130_fd_sc_hs__xnor2_1 _06834_ (.A(net2927),
    .B(net2633),
    .Y(_01407_));
 sky130_fd_sc_hs__nor2_1 _06835_ (.A(net2634),
    .B(_01360_),
    .Y(_01408_));
 sky130_fd_sc_hs__a21oi_2 _06836_ (.A1(net2613),
    .A2(_01407_),
    .B1(_01408_),
    .Y(_01409_));
 sky130_fd_sc_hs__nand2_1 _06837_ (.A(_01406_),
    .B(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hs__inv_1 _06838_ (.A(net2634),
    .Y(_01411_));
 sky130_fd_sc_hs__nand4_1 _06839_ (.A(net3841),
    .B(net2923),
    .C(_01411_),
    .D(net2616),
    .Y(_01412_));
 sky130_fd_sc_hs__nand2_1 _06840_ (.A(_01410_),
    .B(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hs__nand2_2 _06841_ (.A(_01391_),
    .B(_01413_),
    .Y(_01414_));
 sky130_fd_sc_hs__nand3_1 _06842_ (.A(_01387_),
    .B(_01409_),
    .C(_01390_),
    .Y(_01415_));
 sky130_fd_sc_hs__nand2_2 _06843_ (.A(_01414_),
    .B(_01415_),
    .Y(_01416_));
 sky130_fd_sc_hs__nor2_4 _06844_ (.A(_01416_),
    .B(_01405_),
    .Y(_01417_));
 sky130_fd_sc_hs__nand2_2 _06845_ (.A(_01399_),
    .B(_01417_),
    .Y(_01418_));
 sky130_fd_sc_hs__nand2_1 _06846_ (.A(_01361_),
    .B(_01366_),
    .Y(_01419_));
 sky130_fd_sc_hs__nor2_1 _06847_ (.A(_01393_),
    .B(_01419_),
    .Y(_01420_));
 sky130_fd_sc_hs__a21oi_1 _06848_ (.A1(_01420_),
    .A2(net2632),
    .B1(net2597),
    .Y(_01421_));
 sky130_fd_sc_hs__nand4_1 _06849_ (.A(net2599),
    .B(_01403_),
    .C(net2605),
    .D(net2606),
    .Y(_01422_));
 sky130_fd_sc_hs__o21ai_2 _06850_ (.A1(net2606),
    .A2(_01421_),
    .B1(_01422_),
    .Y(_01423_));
 sky130_fd_sc_hs__inv_1 _06851_ (.A(_01423_),
    .Y(_01424_));
 sky130_fd_sc_hs__nand2_2 _06852_ (.A(_01418_),
    .B(_01424_),
    .Y(_01425_));
 sky130_fd_sc_hs__nand2_2 _06853_ (.A(_01425_),
    .B(net2862),
    .Y(_01426_));
 sky130_fd_sc_hs__nand3_2 _06854_ (.A(_01418_),
    .B(net2891),
    .C(_01424_),
    .Y(_01427_));
 sky130_fd_sc_hs__o21ai_1 _06855_ (.A1(net2999),
    .A2(net3043),
    .B1(net2965),
    .Y(_01428_));
 sky130_fd_sc_hs__xnor2_1 _06856_ (.A(net3045),
    .B(_01428_),
    .Y(_01429_));
 sky130_fd_sc_hs__nand2_1 _06857_ (.A(net2563),
    .B(net2568),
    .Y(_01430_));
 sky130_fd_sc_hs__inv_1 _06858_ (.A(_01430_),
    .Y(_01431_));
 sky130_fd_sc_hs__nand4_2 _06859_ (.A(_01426_),
    .B(_01427_),
    .C(net2921),
    .D(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hs__o21ai_2 _06860_ (.A1(net2567),
    .A2(net2545),
    .B1(net2553),
    .Y(_01433_));
 sky130_fd_sc_hs__inv_1 _06861_ (.A(net2552),
    .Y(_01434_));
 sky130_fd_sc_hs__nand2_1 _06862_ (.A(_01433_),
    .B(_01434_),
    .Y(_01435_));
 sky130_fd_sc_hs__nand3_1 _06863_ (.A(net2553),
    .B(net2552),
    .C(net2567),
    .Y(_01436_));
 sky130_fd_sc_hs__nand2_2 _06864_ (.A(_01435_),
    .B(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hs__nor2_1 _06865_ (.A(net2925),
    .B(net2595),
    .Y(_01438_));
 sky130_fd_sc_hs__o21ai_2 _06866_ (.A1(net2588),
    .A2(_01438_),
    .B1(net2569),
    .Y(_01439_));
 sky130_fd_sc_hs__nand3_1 _06867_ (.A(net2577),
    .B(net2594),
    .C(net2596),
    .Y(_01440_));
 sky130_fd_sc_hs__and2_2 _06868_ (.A(_01439_),
    .B(_01440_),
    .X(_01441_));
 sky130_fd_sc_hs__nand3_1 _06869_ (.A(_01392_),
    .B(_01394_),
    .C(net2863),
    .Y(_01442_));
 sky130_fd_sc_hs__nand2_1 _06870_ (.A(_01441_),
    .B(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hs__nand4_1 _06871_ (.A(_01392_),
    .B(_01394_),
    .C(net2863),
    .D(net2594),
    .Y(_01444_));
 sky130_fd_sc_hs__and2_2 _06872_ (.A(_01443_),
    .B(_01444_),
    .X(_01445_));
 sky130_fd_sc_hs__nand2_2 _06873_ (.A(_01425_),
    .B(_01445_),
    .Y(_01446_));
 sky130_fd_sc_hs__inv_1 _06874_ (.A(_01441_),
    .Y(_01447_));
 sky130_fd_sc_hs__nand3_1 _06875_ (.A(_01418_),
    .B(_01447_),
    .C(_01424_),
    .Y(_01448_));
 sky130_fd_sc_hs__nand2_2 _06876_ (.A(_01446_),
    .B(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hs__and2_2 _06877_ (.A(_01437_),
    .B(_01449_),
    .X(_01450_));
 sky130_fd_sc_hs__nand2_2 _06878_ (.A(_01432_),
    .B(_01450_),
    .Y(_01451_));
 sky130_fd_sc_hs__nand2_1 _06879_ (.A(net2553),
    .B(_01434_),
    .Y(_01452_));
 sky130_fd_sc_hs__o21ai_1 _06880_ (.A1(_01424_),
    .A2(_01452_),
    .B1(net2562),
    .Y(_01453_));
 sky130_fd_sc_hs__nand2_2 _06881_ (.A(_01453_),
    .B(net2533),
    .Y(_01454_));
 sky130_fd_sc_hs__nand2_2 _06882_ (.A(_01454_),
    .B(_01451_),
    .Y(_01455_));
 sky130_fd_sc_hs__nand2_2 _06883_ (.A(_01455_),
    .B(net2922),
    .Y(_01456_));
 sky130_fd_sc_hs__inv_1 _06884_ (.A(net2922),
    .Y(_01457_));
 sky130_fd_sc_hs__nand3_1 _06885_ (.A(_01451_),
    .B(_01457_),
    .C(_01454_),
    .Y(_01458_));
 sky130_fd_sc_hs__o31ai_1 _06886_ (.A1(net3133),
    .A2(net3140),
    .A3(net2994),
    .B1(net2965),
    .Y(_01459_));
 sky130_fd_sc_hs__xnor2_1 _06887_ (.A(net3047),
    .B(_01459_),
    .Y(_01460_));
 sky130_fd_sc_hs__and2_2 _06888_ (.A(_01426_),
    .B(net2527),
    .X(_01461_));
 sky130_fd_sc_hs__nand4_2 _06889_ (.A(_01456_),
    .B(_01458_),
    .C(net2920),
    .D(net2510),
    .Y(_01462_));
 sky130_fd_sc_hs__xnor2_1 _06890_ (.A(net2891),
    .B(_01430_),
    .Y(_01463_));
 sky130_fd_sc_hs__nand2_1 _06891_ (.A(net3840),
    .B(_01463_),
    .Y(_01464_));
 sky130_fd_sc_hs__o21ai_2 _06892_ (.A1(net2544),
    .A2(net3839),
    .B1(_01464_),
    .Y(_01465_));
 sky130_fd_sc_hs__nand3_1 _06893_ (.A(_01465_),
    .B(_01461_),
    .C(net2922),
    .Y(_01466_));
 sky130_fd_sc_hs__o21a_1 _06894_ (.A1(_01431_),
    .A2(net3839),
    .B1(_01464_),
    .X(_01467_));
 sky130_fd_sc_hs__nand3_1 _06895_ (.A(_01426_),
    .B(net2527),
    .C(net2921),
    .Y(_01468_));
 sky130_fd_sc_hs__nand2_1 _06896_ (.A(_01467_),
    .B(_01468_),
    .Y(_01469_));
 sky130_fd_sc_hs__nand2_1 _06897_ (.A(_01466_),
    .B(_01469_),
    .Y(_01470_));
 sky130_fd_sc_hs__nand2_2 _06898_ (.A(_01455_),
    .B(_01470_),
    .Y(_01471_));
 sky130_fd_sc_hs__nand3_1 _06899_ (.A(_01451_),
    .B(_01467_),
    .C(_01454_),
    .Y(_01472_));
 sky130_fd_sc_hs__nand2_2 _06900_ (.A(_01471_),
    .B(_01472_),
    .Y(_01473_));
 sky130_fd_sc_hs__nor2_2 _06901_ (.A(net2551),
    .B(_01468_),
    .Y(_01474_));
 sky130_fd_sc_hs__inv_1 _06902_ (.A(net2511),
    .Y(_01475_));
 sky130_fd_sc_hs__nand2_1 _06903_ (.A(_01474_),
    .B(_01475_),
    .Y(_01476_));
 sky130_fd_sc_hs__nand2_1 _06904_ (.A(net2512),
    .B(net2511),
    .Y(_01477_));
 sky130_fd_sc_hs__nand2_1 _06905_ (.A(_01476_),
    .B(_01477_),
    .Y(_01478_));
 sky130_fd_sc_hs__nand2_1 _06906_ (.A(_01478_),
    .B(_01455_),
    .Y(_01479_));
 sky130_fd_sc_hs__nand3_1 _06907_ (.A(net2491),
    .B(_01475_),
    .C(net2519),
    .Y(_01480_));
 sky130_fd_sc_hs__nand2_2 _06908_ (.A(_01479_),
    .B(_01480_),
    .Y(_01481_));
 sky130_fd_sc_hs__nor2_4 _06909_ (.A(_01473_),
    .B(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hs__nand2_2 _06910_ (.A(_01462_),
    .B(_01482_),
    .Y(_01483_));
 sky130_fd_sc_hs__inv_1 _06911_ (.A(net2520),
    .Y(_01484_));
 sky130_fd_sc_hs__nand3b_1 _06912_ (.A_N(_01477_),
    .B(net2487),
    .C(_01484_),
    .Y(_01485_));
 sky130_fd_sc_hs__nand2_1 _06913_ (.A(net2501),
    .B(net2520),
    .Y(_01486_));
 sky130_fd_sc_hs__nand2_2 _06914_ (.A(_01485_),
    .B(_01486_),
    .Y(_01487_));
 sky130_fd_sc_hs__inv_2 _06915_ (.A(_01487_),
    .Y(_01488_));
 sky130_fd_sc_hs__nand2_2 _06916_ (.A(_01488_),
    .B(_01483_),
    .Y(_01489_));
 sky130_fd_sc_hs__nand2_2 _06917_ (.A(net2920),
    .B(_01489_),
    .Y(_01490_));
 sky130_fd_sc_hs__inv_1 _06918_ (.A(net2920),
    .Y(_01491_));
 sky130_fd_sc_hs__nand3_2 _06919_ (.A(_01483_),
    .B(_01491_),
    .C(_01488_),
    .Y(_01492_));
 sky130_fd_sc_hs__and2_1 _06920_ (.A(net2966),
    .B(net3043),
    .X(_01493_));
 sky130_fd_sc_hs__xnor2_1 _06921_ (.A(net3133),
    .B(_01493_),
    .Y(_01494_));
 sky130_fd_sc_hs__and2_2 _06922_ (.A(net2480),
    .B(net2486),
    .X(_01495_));
 sky130_fd_sc_hs__nand4_2 _06923_ (.A(_01490_),
    .B(_01492_),
    .C(_01494_),
    .D(net2464),
    .Y(_01496_));
 sky130_fd_sc_hs__inv_1 _06924_ (.A(net2466),
    .Y(_01497_));
 sky130_fd_sc_hs__and2_1 _06925_ (.A(net2467),
    .B(_01497_),
    .X(_01498_));
 sky130_fd_sc_hs__nand2_2 _06926_ (.A(_01489_),
    .B(_01498_),
    .Y(_01499_));
 sky130_fd_sc_hs__nand2_2 _06927_ (.A(_01499_),
    .B(net2465),
    .Y(_01500_));
 sky130_fd_sc_hs__and2_2 _06928_ (.A(net2422),
    .B(net2447),
    .X(_01501_));
 sky130_fd_sc_hs__o21ai_2 _06929_ (.A1(_01487_),
    .A2(_01482_),
    .B1(net2468),
    .Y(_01502_));
 sky130_fd_sc_hs__nand2_1 _06930_ (.A(_01502_),
    .B(net2466),
    .Y(_01503_));
 sky130_fd_sc_hs__nand2_2 _06931_ (.A(_01499_),
    .B(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hs__nand2_1 _06932_ (.A(_01495_),
    .B(net2920),
    .Y(_01505_));
 sky130_fd_sc_hs__inv_1 _06933_ (.A(net2510),
    .Y(_01506_));
 sky130_fd_sc_hs__nand2_1 _06934_ (.A(net2479),
    .B(_01506_),
    .Y(_01507_));
 sky130_fd_sc_hs__nand3_1 _06935_ (.A(net3795),
    .B(net2922),
    .C(net2510),
    .Y(_01508_));
 sky130_fd_sc_hs__and2_2 _06936_ (.A(_01507_),
    .B(_01508_),
    .X(_01509_));
 sky130_fd_sc_hs__nand2_1 _06937_ (.A(_01505_),
    .B(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hs__nand4_1 _06938_ (.A(net2480),
    .B(net2486),
    .C(net2920),
    .D(net2500),
    .Y(_01511_));
 sky130_fd_sc_hs__nand2_1 _06939_ (.A(_01510_),
    .B(_01511_),
    .Y(_01512_));
 sky130_fd_sc_hs__nand2_2 _06940_ (.A(_01489_),
    .B(_01512_),
    .Y(_01513_));
 sky130_fd_sc_hs__nand3_1 _06941_ (.A(_01483_),
    .B(_01488_),
    .C(_01509_),
    .Y(_01514_));
 sky130_fd_sc_hs__and2_2 _06942_ (.A(_01513_),
    .B(_01514_),
    .X(_01515_));
 sky130_fd_sc_hs__nand4_1 _06943_ (.A(net2423),
    .B(_01501_),
    .C(net2421),
    .D(_01515_),
    .Y(_01516_));
 sky130_fd_sc_hs__nand2_1 _06944_ (.A(net2423),
    .B(_01515_),
    .Y(_01517_));
 sky130_fd_sc_hs__and2_1 _06945_ (.A(net2438),
    .B(net2430),
    .X(_01518_));
 sky130_fd_sc_hs__nand2_1 _06946_ (.A(_01517_),
    .B(_01518_),
    .Y(_01519_));
 sky130_fd_sc_hs__nand2_2 _06947_ (.A(_01516_),
    .B(_01519_),
    .Y(_01520_));
 sky130_fd_sc_hs__nand2_2 _06948_ (.A(_01513_),
    .B(_01514_),
    .Y(_01521_));
 sky130_fd_sc_hs__nor2_4 _06949_ (.A(_01504_),
    .B(_01521_),
    .Y(_01522_));
 sky130_fd_sc_hs__nand2_2 _06950_ (.A(_01522_),
    .B(_01496_),
    .Y(_01523_));
 sky130_fd_sc_hs__nand2_2 _06951_ (.A(_01500_),
    .B(net2447),
    .Y(_01524_));
 sky130_fd_sc_hs__nand2_2 _06952_ (.A(_01523_),
    .B(net2408),
    .Y(_01525_));
 sky130_fd_sc_hs__inv_1 _06953_ (.A(net2464),
    .Y(_01526_));
 sky130_fd_sc_hs__nand2_1 _06954_ (.A(net2431),
    .B(_01526_),
    .Y(_01527_));
 sky130_fd_sc_hs__nand3_1 _06955_ (.A(net4866),
    .B(net2920),
    .C(net2464),
    .Y(_01528_));
 sky130_fd_sc_hs__and2_1 _06956_ (.A(_01527_),
    .B(_01528_),
    .X(_01529_));
 sky130_fd_sc_hs__and2_2 _06957_ (.A(_01490_),
    .B(_01492_),
    .X(_01530_));
 sky130_fd_sc_hs__nand2_1 _06958_ (.A(_01530_),
    .B(_01494_),
    .Y(_01531_));
 sky130_fd_sc_hs__nand2_1 _06959_ (.A(_01529_),
    .B(_01531_),
    .Y(_01532_));
 sky130_fd_sc_hs__nand4_1 _06960_ (.A(net2431),
    .B(net2439),
    .C(net2919),
    .D(_01526_),
    .Y(_01533_));
 sky130_fd_sc_hs__nand2_1 _06961_ (.A(_01532_),
    .B(_01533_),
    .Y(_01534_));
 sky130_fd_sc_hs__nand2_2 _06962_ (.A(_01525_),
    .B(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hs__nand3_1 _06963_ (.A(_01523_),
    .B(net2408),
    .C(_01529_),
    .Y(_01536_));
 sky130_fd_sc_hs__nand2_2 _06964_ (.A(_01535_),
    .B(_01536_),
    .Y(_01537_));
 sky130_fd_sc_hs__inv_1 _06965_ (.A(_01494_),
    .Y(_01538_));
 sky130_fd_sc_hs__nand3_1 _06966_ (.A(net4927),
    .B(_01492_),
    .C(net2464),
    .Y(_01539_));
 sky130_fd_sc_hs__nor2_1 _06967_ (.A(_01538_),
    .B(_01539_),
    .Y(_01540_));
 sky130_fd_sc_hs__nand2_1 _06968_ (.A(_01540_),
    .B(net2418),
    .Y(_01541_));
 sky130_fd_sc_hs__nand2_1 _06969_ (.A(_01541_),
    .B(_01517_),
    .Y(_01542_));
 sky130_fd_sc_hs__nand2_2 _06970_ (.A(_01542_),
    .B(_01525_),
    .Y(_01543_));
 sky130_fd_sc_hs__nand3_1 _06971_ (.A(net2398),
    .B(net2408),
    .C(net2418),
    .Y(_01544_));
 sky130_fd_sc_hs__nand2_2 _06972_ (.A(_01543_),
    .B(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hs__nor2_4 _06973_ (.A(_01537_),
    .B(_01545_),
    .Y(_01546_));
 sky130_fd_sc_hs__nand2_2 _06974_ (.A(_01525_),
    .B(_01494_),
    .Y(_01547_));
 sky130_fd_sc_hs__o211ai_2 _06975_ (.A1(_01521_),
    .A2(net4920),
    .B1(_01538_),
    .C1(_01524_),
    .Y(_01548_));
 sky130_fd_sc_hs__nand2_1 _06976_ (.A(net2966),
    .B(net2994),
    .Y(_01549_));
 sky130_fd_sc_hs__xnor2_1 _06977_ (.A(net3140),
    .B(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hs__clkinv_1 _06978_ (.A(_01550_),
    .Y(_01551_));
 sky130_fd_sc_hs__nand4_2 _06979_ (.A(_01547_),
    .B(_01548_),
    .C(_01551_),
    .D(net2417),
    .Y(_01552_));
 sky130_fd_sc_hs__o21ai_1 _06980_ (.A1(_01520_),
    .A2(_01546_),
    .B1(net3800),
    .Y(_01553_));
 sky130_fd_sc_hs__nand2_1 _06981_ (.A(_01553_),
    .B(net2370),
    .Y(_01554_));
 sky130_fd_sc_hs__nand2_1 _06982_ (.A(_01518_),
    .B(net2420),
    .Y(_01555_));
 sky130_fd_sc_hs__a21oi_1 _06983_ (.A1(_01555_),
    .A2(net2408),
    .B1(net2406),
    .Y(_01556_));
 sky130_fd_sc_hs__nand2_1 _06984_ (.A(_01556_),
    .B(net2418),
    .Y(_01557_));
 sky130_fd_sc_hs__o21ai_1 _06985_ (.A1(_01501_),
    .A2(net2410),
    .B1(net2423),
    .Y(_01558_));
 sky130_fd_sc_hs__nand2_1 _06986_ (.A(_01558_),
    .B(net2419),
    .Y(_01559_));
 sky130_fd_sc_hs__nand2_1 _06987_ (.A(_01557_),
    .B(_01559_),
    .Y(_01560_));
 sky130_fd_sc_hs__and2_2 _06988_ (.A(_01535_),
    .B(_01536_),
    .X(_01561_));
 sky130_fd_sc_hs__o211ai_1 _06989_ (.A1(_01520_),
    .A2(_01560_),
    .B1(_01561_),
    .C1(net2368),
    .Y(_01562_));
 sky130_fd_sc_hs__nand2_1 _06990_ (.A(_01554_),
    .B(_01562_),
    .Y(_01563_));
 sky130_fd_sc_hs__nand2_2 _06991_ (.A(_01552_),
    .B(_01546_),
    .Y(_01564_));
 sky130_fd_sc_hs__inv_1 _06992_ (.A(_01520_),
    .Y(_01565_));
 sky130_fd_sc_hs__nand2_2 _06993_ (.A(_01564_),
    .B(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hs__inv_2 _06994_ (.A(net2417),
    .Y(_01567_));
 sky130_fd_sc_hs__nand2_1 _06995_ (.A(_01567_),
    .B(_01538_),
    .Y(_01568_));
 sky130_fd_sc_hs__nand2_1 _06996_ (.A(_01568_),
    .B(net2407),
    .Y(_01569_));
 sky130_fd_sc_hs__nand2_1 _06997_ (.A(net2389),
    .B(_01569_),
    .Y(_01570_));
 sky130_fd_sc_hs__nand3_1 _06998_ (.A(net2397),
    .B(_01567_),
    .C(net2409),
    .Y(_01571_));
 sky130_fd_sc_hs__nand2_2 _06999_ (.A(_01570_),
    .B(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hs__nand3_2 _07000_ (.A(_01547_),
    .B(_01551_),
    .C(net2396),
    .Y(_01573_));
 sky130_fd_sc_hs__xnor2_2 _07001_ (.A(_01572_),
    .B(_01573_),
    .Y(_01574_));
 sky130_fd_sc_hs__nand2_1 _07002_ (.A(_01560_),
    .B(_01561_),
    .Y(_01575_));
 sky130_fd_sc_hs__nand3_1 _07003_ (.A(_01575_),
    .B(_01572_),
    .C(_01565_),
    .Y(_01576_));
 sky130_fd_sc_hs__a21boi_2 _07004_ (.A1(_01566_),
    .A2(_01574_),
    .B1_N(_01576_),
    .Y(_01577_));
 sky130_fd_sc_hs__nor2_2 _07005_ (.A(_01563_),
    .B(_01577_),
    .Y(_01578_));
 sky130_fd_sc_hs__nand3_2 _07006_ (.A(_01564_),
    .B(_01551_),
    .C(_01565_),
    .Y(_01579_));
 sky130_fd_sc_hs__o21ai_2 _07007_ (.A1(_01520_),
    .A2(_01546_),
    .B1(_01550_),
    .Y(_01580_));
 sky130_fd_sc_hs__nand2_2 _07008_ (.A(_01579_),
    .B(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hs__nor2_1 _07009_ (.A(net3233),
    .B(net3144),
    .Y(_01582_));
 sky130_fd_sc_hs__nand4_1 _07010_ (.A(_01582_),
    .B(net3231),
    .C(net3229),
    .D(net3189),
    .Y(_01583_));
 sky130_fd_sc_hs__inv_1 _07011_ (.A(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hs__a31o_1 _07012_ (.A1(_01584_),
    .A2(net3094),
    .A3(net3093),
    .B1(net2944),
    .X(_01585_));
 sky130_fd_sc_hs__xnor2_1 _07013_ (.A(net3134),
    .B(_01585_),
    .Y(_01586_));
 sky130_fd_sc_hs__nand2_1 _07014_ (.A(net2381),
    .B(net2396),
    .Y(_01587_));
 sky130_fd_sc_hs__inv_1 _07015_ (.A(_01587_),
    .Y(_01588_));
 sky130_fd_sc_hs__nand3_2 _07016_ (.A(_01581_),
    .B(_01586_),
    .C(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hs__nand2_2 _07017_ (.A(_01589_),
    .B(_01578_),
    .Y(_01590_));
 sky130_fd_sc_hs__inv_1 _07018_ (.A(net2313),
    .Y(_01591_));
 sky130_fd_sc_hs__inv_1 _07019_ (.A(net3798),
    .Y(_01592_));
 sky130_fd_sc_hs__nand2_1 _07020_ (.A(_01562_),
    .B(net2369),
    .Y(_01593_));
 sky130_fd_sc_hs__and2_2 _07021_ (.A(_01593_),
    .B(net2352),
    .X(_01594_));
 sky130_fd_sc_hs__and2_1 _07022_ (.A(_01554_),
    .B(_01562_),
    .X(_01595_));
 sky130_fd_sc_hs__a31oi_1 _07023_ (.A1(_01592_),
    .A2(net2322),
    .A3(net2344),
    .B1(_01595_),
    .Y(_01596_));
 sky130_fd_sc_hs__nor2_1 _07024_ (.A(_01591_),
    .B(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hs__inv_2 _07025_ (.A(_01597_),
    .Y(_01598_));
 sky130_fd_sc_hs__inv_2 _07026_ (.A(_01594_),
    .Y(_01599_));
 sky130_fd_sc_hs__nand2_2 _07027_ (.A(_01590_),
    .B(_01599_),
    .Y(_01600_));
 sky130_fd_sc_hs__nand2_2 _07028_ (.A(_01600_),
    .B(_01586_),
    .Y(_01601_));
 sky130_fd_sc_hs__inv_1 _07029_ (.A(_01586_),
    .Y(_01602_));
 sky130_fd_sc_hs__nand3_2 _07030_ (.A(_01590_),
    .B(_01602_),
    .C(_01599_),
    .Y(_01603_));
 sky130_fd_sc_hs__nand2_1 _07031_ (.A(net2966),
    .B(net3034),
    .Y(_01604_));
 sky130_fd_sc_hs__xnor2_1 _07032_ (.A(net3135),
    .B(_01604_),
    .Y(_01605_));
 sky130_fd_sc_hs__nand4_2 _07033_ (.A(_01601_),
    .B(_01603_),
    .C(_01605_),
    .D(net2333),
    .Y(_01606_));
 sky130_fd_sc_hs__nand2_1 _07034_ (.A(_01566_),
    .B(_01551_),
    .Y(_01607_));
 sky130_fd_sc_hs__nand2_1 _07035_ (.A(_01607_),
    .B(net2366),
    .Y(_01608_));
 sky130_fd_sc_hs__inv_1 _07036_ (.A(net2367),
    .Y(_01609_));
 sky130_fd_sc_hs__nand2_1 _07037_ (.A(net2345),
    .B(_01609_),
    .Y(_01610_));
 sky130_fd_sc_hs__and2_2 _07038_ (.A(_01608_),
    .B(_01610_),
    .X(_01611_));
 sky130_fd_sc_hs__nand2_1 _07039_ (.A(_01581_),
    .B(_01586_),
    .Y(_01612_));
 sky130_fd_sc_hs__nand2_1 _07040_ (.A(_01611_),
    .B(_01612_),
    .Y(_01613_));
 sky130_fd_sc_hs__and2_1 _07041_ (.A(_01579_),
    .B(_01580_),
    .X(_01614_));
 sky130_fd_sc_hs__nor2_1 _07042_ (.A(_01602_),
    .B(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hs__nand2_1 _07043_ (.A(_01608_),
    .B(_01610_),
    .Y(_01616_));
 sky130_fd_sc_hs__nand2_1 _07044_ (.A(_01615_),
    .B(_01616_),
    .Y(_01617_));
 sky130_fd_sc_hs__nand2_1 _07045_ (.A(_01613_),
    .B(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hs__nand2_1 _07046_ (.A(_01600_),
    .B(_01618_),
    .Y(_01619_));
 sky130_fd_sc_hs__nand3_1 _07047_ (.A(_01590_),
    .B(net2312),
    .C(_01599_),
    .Y(_01620_));
 sky130_fd_sc_hs__nand2_2 _07048_ (.A(_01619_),
    .B(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hs__inv_1 _07049_ (.A(net2285),
    .Y(_01622_));
 sky130_fd_sc_hs__nand2_1 _07050_ (.A(net2293),
    .B(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hs__o211ai_1 _07051_ (.A1(_01595_),
    .A2(_01594_),
    .B1(_01592_),
    .C1(net2322),
    .Y(_01624_));
 sky130_fd_sc_hs__a21o_1 _07052_ (.A1(net2322),
    .A2(net2344),
    .B1(_01592_),
    .X(_01625_));
 sky130_fd_sc_hs__nand2_1 _07053_ (.A(_01624_),
    .B(_01625_),
    .Y(_01626_));
 sky130_fd_sc_hs__o21ai_1 _07054_ (.A1(_01598_),
    .A2(_01623_),
    .B1(net2306),
    .Y(_01627_));
 sky130_fd_sc_hs__nor2_4 _07055_ (.A(_01626_),
    .B(_01621_),
    .Y(_01628_));
 sky130_fd_sc_hs__nand2_2 _07056_ (.A(_01628_),
    .B(_01606_),
    .Y(_01629_));
 sky130_fd_sc_hs__and2_1 _07057_ (.A(_01627_),
    .B(_01629_),
    .X(_01630_));
 sky130_fd_sc_hs__inv_2 _07058_ (.A(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hs__nand2_2 _07059_ (.A(_01598_),
    .B(_01629_),
    .Y(_01632_));
 sky130_fd_sc_hs__nand2_2 _07060_ (.A(_01632_),
    .B(_01605_),
    .Y(_01633_));
 sky130_fd_sc_hs__inv_1 _07061_ (.A(_01605_),
    .Y(_01634_));
 sky130_fd_sc_hs__nand3_2 _07062_ (.A(_01598_),
    .B(_01634_),
    .C(_01629_),
    .Y(_01635_));
 sky130_fd_sc_hs__inv_1 _07063_ (.A(net3138),
    .Y(_01636_));
 sky130_fd_sc_hs__o31ai_1 _07064_ (.A1(net3142),
    .A2(net3141),
    .A3(_01583_),
    .B1(net2966),
    .Y(_01637_));
 sky130_fd_sc_hs__xnor2_1 _07065_ (.A(_01636_),
    .B(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hs__nand2_1 _07066_ (.A(_01601_),
    .B(_01603_),
    .Y(_01639_));
 sky130_fd_sc_hs__clkdlyinv3sd1_1 _07067_ (.A(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hs__nand4_4 _07068_ (.A(_01633_),
    .B(_01635_),
    .C(net2918),
    .D(_01640_),
    .Y(_01641_));
 sky130_fd_sc_hs__xnor2_1 _07069_ (.A(_01586_),
    .B(net2333),
    .Y(_01642_));
 sky130_fd_sc_hs__nand2_1 _07070_ (.A(net4896),
    .B(_01642_),
    .Y(_01643_));
 sky130_fd_sc_hs__o21ai_2 _07071_ (.A1(net2333),
    .A2(_01600_),
    .B1(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hs__nand3_2 _07072_ (.A(net2299),
    .B(net2307),
    .C(_01605_),
    .Y(_01645_));
 sky130_fd_sc_hs__xnor2_2 _07073_ (.A(_01645_),
    .B(_01644_),
    .Y(_01646_));
 sky130_fd_sc_hs__nand2_1 _07074_ (.A(_01632_),
    .B(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hs__nand3_2 _07075_ (.A(_01629_),
    .B(_01644_),
    .C(_01598_),
    .Y(_01648_));
 sky130_fd_sc_hs__nand2_2 _07076_ (.A(_01647_),
    .B(_01648_),
    .Y(_01649_));
 sky130_fd_sc_hs__nand2_1 _07077_ (.A(net3832),
    .B(net2251),
    .Y(_01650_));
 sky130_fd_sc_hs__o21ai_1 _07078_ (.A1(_01597_),
    .A2(_01628_),
    .B1(_01606_),
    .Y(_01651_));
 sky130_fd_sc_hs__nand2_1 _07079_ (.A(_01651_),
    .B(_01622_),
    .Y(_01652_));
 sky130_fd_sc_hs__nand3_1 _07080_ (.A(net2293),
    .B(net2285),
    .C(net2300),
    .Y(_01653_));
 sky130_fd_sc_hs__nand2_1 _07081_ (.A(_01652_),
    .B(_01653_),
    .Y(_01654_));
 sky130_fd_sc_hs__o21bai_1 _07082_ (.A1(_01631_),
    .A2(_01650_),
    .B1_N(net2256),
    .Y(_01655_));
 sky130_fd_sc_hs__and2_2 _07083_ (.A(_01649_),
    .B(_01654_),
    .X(_01656_));
 sky130_fd_sc_hs__nand2_2 _07084_ (.A(_01656_),
    .B(_01641_),
    .Y(_01657_));
 sky130_fd_sc_hs__and2_2 _07085_ (.A(_01655_),
    .B(net2232),
    .X(_01658_));
 sky130_fd_sc_hs__o21ai_1 _07086_ (.A1(_01630_),
    .A2(net2238),
    .B1(net2252),
    .Y(_01659_));
 sky130_fd_sc_hs__inv_1 _07087_ (.A(net2251),
    .Y(_01660_));
 sky130_fd_sc_hs__nand2_1 _07088_ (.A(_01660_),
    .B(_01659_),
    .Y(_01661_));
 sky130_fd_sc_hs__o211ai_1 _07089_ (.A1(net2256),
    .A2(_01630_),
    .B1(net2251),
    .C1(net2252),
    .Y(_01662_));
 sky130_fd_sc_hs__nand2_1 _07090_ (.A(_01661_),
    .B(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hs__xnor2_1 _07091_ (.A(_01640_),
    .B(_01633_),
    .Y(_01664_));
 sky130_fd_sc_hs__and2_1 _07092_ (.A(_01633_),
    .B(net4929),
    .X(_01665_));
 sky130_fd_sc_hs__nand2_1 _07093_ (.A(_01665_),
    .B(net2918),
    .Y(_01666_));
 sky130_fd_sc_hs__nand2_1 _07094_ (.A(_01664_),
    .B(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hs__nand4_1 _07095_ (.A(net2257),
    .B(net2266),
    .C(net2918),
    .D(net2292),
    .Y(_01668_));
 sky130_fd_sc_hs__nand2_1 _07096_ (.A(_01667_),
    .B(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hs__nand2_2 _07097_ (.A(_01657_),
    .B(_01631_),
    .Y(_01670_));
 sky130_fd_sc_hs__nand2_2 _07098_ (.A(_01669_),
    .B(_01670_),
    .Y(_01671_));
 sky130_fd_sc_hs__nand3_1 _07099_ (.A(_01657_),
    .B(_01631_),
    .C(net2250),
    .Y(_01672_));
 sky130_fd_sc_hs__nand2_2 _07100_ (.A(_01671_),
    .B(_01672_),
    .Y(_01673_));
 sky130_fd_sc_hs__nor2_4 _07101_ (.A(_01673_),
    .B(_01663_),
    .Y(_01674_));
 sky130_fd_sc_hs__nand2_2 _07102_ (.A(_01670_),
    .B(net2918),
    .Y(_01675_));
 sky130_fd_sc_hs__inv_1 _07103_ (.A(net2918),
    .Y(_01676_));
 sky130_fd_sc_hs__nand3_2 _07104_ (.A(_01657_),
    .B(_01676_),
    .C(_01631_),
    .Y(_01677_));
 sky130_fd_sc_hs__nor2_1 _07105_ (.A(net3032),
    .B(net2944),
    .Y(_01678_));
 sky130_fd_sc_hs__xnor2_1 _07106_ (.A(net3141),
    .B(_01678_),
    .Y(_01679_));
 sky130_fd_sc_hs__nand4_2 _07107_ (.A(_01675_),
    .B(_01677_),
    .C(net2890),
    .D(net2249),
    .Y(_01680_));
 sky130_fd_sc_hs__o21ai_1 _07108_ (.A1(_01658_),
    .A2(_01674_),
    .B1(_01680_),
    .Y(_01681_));
 sky130_fd_sc_hs__nand2_1 _07109_ (.A(_01681_),
    .B(net2207),
    .Y(_01682_));
 sky130_fd_sc_hs__and2_1 _07110_ (.A(_01661_),
    .B(_01662_),
    .X(_01683_));
 sky130_fd_sc_hs__and2_2 _07111_ (.A(_01671_),
    .B(_01672_),
    .X(_01684_));
 sky130_fd_sc_hs__o211ai_1 _07112_ (.A1(_01683_),
    .A2(_01658_),
    .B1(_01684_),
    .C1(_01680_),
    .Y(_01685_));
 sky130_fd_sc_hs__nand2_1 _07113_ (.A(_01682_),
    .B(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hs__nand2_2 _07114_ (.A(_01680_),
    .B(_01674_),
    .Y(_01687_));
 sky130_fd_sc_hs__inv_1 _07115_ (.A(_01658_),
    .Y(_01688_));
 sky130_fd_sc_hs__nand2_2 _07116_ (.A(_01687_),
    .B(_01688_),
    .Y(_01689_));
 sky130_fd_sc_hs__nand2_1 _07117_ (.A(net4871),
    .B(_01635_),
    .Y(_01690_));
 sky130_fd_sc_hs__xnor2_1 _07118_ (.A(_01676_),
    .B(_01690_),
    .Y(_01691_));
 sky130_fd_sc_hs__nand2_1 _07119_ (.A(net4904),
    .B(_01691_),
    .Y(_01692_));
 sky130_fd_sc_hs__nand3_1 _07120_ (.A(net3804),
    .B(_01631_),
    .C(_01690_),
    .Y(_01693_));
 sky130_fd_sc_hs__and2_4 _07121_ (.A(_01692_),
    .B(_01693_),
    .X(_01694_));
 sky130_fd_sc_hs__nand3_1 _07122_ (.A(_01675_),
    .B(_01677_),
    .C(net2890),
    .Y(_01695_));
 sky130_fd_sc_hs__nor2_1 _07123_ (.A(_01694_),
    .B(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hs__and2_1 _07124_ (.A(_01695_),
    .B(_01694_),
    .X(_01697_));
 sky130_fd_sc_hs__nor2_2 _07125_ (.A(_01696_),
    .B(_01697_),
    .Y(_01698_));
 sky130_fd_sc_hs__nand2_1 _07126_ (.A(_01689_),
    .B(_01698_),
    .Y(_01699_));
 sky130_fd_sc_hs__nand2_1 _07127_ (.A(_01684_),
    .B(_01683_),
    .Y(_01700_));
 sky130_fd_sc_hs__nand3b_1 _07128_ (.A_N(net2206),
    .B(_01688_),
    .C(_01700_),
    .Y(_01701_));
 sky130_fd_sc_hs__and2_2 _07129_ (.A(_01701_),
    .B(_01699_),
    .X(_01702_));
 sky130_fd_sc_hs__nor2_4 _07130_ (.A(_01686_),
    .B(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hs__nand2_2 _07131_ (.A(_01689_),
    .B(net2890),
    .Y(_01704_));
 sky130_fd_sc_hs__nor2_1 _07132_ (.A(_01584_),
    .B(net2945),
    .Y(_01705_));
 sky130_fd_sc_hs__xnor2_1 _07133_ (.A(net3142),
    .B(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hs__nand2_1 _07134_ (.A(net2217),
    .B(net2227),
    .Y(_01707_));
 sky130_fd_sc_hs__inv_1 _07135_ (.A(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hs__nand3b_1 _07136_ (.A_N(net2890),
    .B(_01688_),
    .C(_01700_),
    .Y(_01709_));
 sky130_fd_sc_hs__nand4_2 _07137_ (.A(_01704_),
    .B(net2889),
    .C(_01708_),
    .D(_01709_),
    .Y(_01710_));
 sky130_fd_sc_hs__nand2_2 _07138_ (.A(_01703_),
    .B(_01710_),
    .Y(_01711_));
 sky130_fd_sc_hs__nand2_1 _07139_ (.A(_01685_),
    .B(net2218),
    .Y(_01712_));
 sky130_fd_sc_hs__and2_1 _07140_ (.A(_01712_),
    .B(_01687_),
    .X(_01713_));
 sky130_fd_sc_hs__inv_1 _07141_ (.A(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hs__nand2_2 _07142_ (.A(_01711_),
    .B(_01714_),
    .Y(_01715_));
 sky130_fd_sc_hs__nand2_2 _07143_ (.A(_01715_),
    .B(net2889),
    .Y(_01716_));
 sky130_fd_sc_hs__inv_1 _07144_ (.A(net2889),
    .Y(_01717_));
 sky130_fd_sc_hs__nand3_1 _07145_ (.A(_01711_),
    .B(_01717_),
    .C(_01714_),
    .Y(_01718_));
 sky130_fd_sc_hs__nor2_1 _07146_ (.A(_01145_),
    .B(net2945),
    .Y(_01719_));
 sky130_fd_sc_hs__xnor2_1 _07147_ (.A(net3144),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hs__and2_2 _07148_ (.A(_01704_),
    .B(net2195),
    .X(_01721_));
 sky130_fd_sc_hs__nand4_1 _07149_ (.A(_01716_),
    .B(_01718_),
    .C(_01720_),
    .D(net2166),
    .Y(_01722_));
 sky130_fd_sc_hs__nand2_1 _07150_ (.A(net2179),
    .B(net2205),
    .Y(_01723_));
 sky130_fd_sc_hs__nand3_1 _07151_ (.A(net2190),
    .B(net2890),
    .C(_01708_),
    .Y(_01724_));
 sky130_fd_sc_hs__and2_2 _07152_ (.A(_01723_),
    .B(_01724_),
    .X(_01725_));
 sky130_fd_sc_hs__nand2_1 _07153_ (.A(_01721_),
    .B(net2889),
    .Y(_01726_));
 sky130_fd_sc_hs__nand2_1 _07154_ (.A(_01725_),
    .B(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hs__nand4_1 _07155_ (.A(_01704_),
    .B(net2889),
    .C(net2205),
    .D(net2196),
    .Y(_01728_));
 sky130_fd_sc_hs__nand2_1 _07156_ (.A(_01727_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hs__nand2_1 _07157_ (.A(_01715_),
    .B(_01729_),
    .Y(_01730_));
 sky130_fd_sc_hs__nand3_1 _07158_ (.A(_01711_),
    .B(net2178),
    .C(_01725_),
    .Y(_01731_));
 sky130_fd_sc_hs__nand2_2 _07159_ (.A(_01730_),
    .B(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hs__o21ai_1 _07160_ (.A1(net2189),
    .A2(_01703_),
    .B1(net2167),
    .Y(_01733_));
 sky130_fd_sc_hs__nand2_1 _07161_ (.A(_01733_),
    .B(net2168),
    .Y(_01734_));
 sky130_fd_sc_hs__inv_1 _07162_ (.A(net2168),
    .Y(_01735_));
 sky130_fd_sc_hs__and2_1 _07163_ (.A(_01735_),
    .B(_01710_),
    .X(_01736_));
 sky130_fd_sc_hs__nand2_2 _07164_ (.A(_01715_),
    .B(_01736_),
    .Y(_01737_));
 sky130_fd_sc_hs__nand2_2 _07165_ (.A(_01737_),
    .B(_01734_),
    .Y(_01738_));
 sky130_fd_sc_hs__nor2_2 _07166_ (.A(_01732_),
    .B(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hs__nand2_2 _07167_ (.A(_01722_),
    .B(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hs__xnor2_4 _07168_ (.A(_01737_),
    .B(net2180),
    .Y(_01741_));
 sky130_fd_sc_hs__nand2_2 _07169_ (.A(_01741_),
    .B(_01740_),
    .Y(_01742_));
 sky130_fd_sc_hs__nand2_2 _07170_ (.A(_01742_),
    .B(_01720_),
    .Y(_01743_));
 sky130_fd_sc_hs__inv_1 _07171_ (.A(_01720_),
    .Y(_01744_));
 sky130_fd_sc_hs__nand3_2 _07172_ (.A(_01744_),
    .B(_01740_),
    .C(_01741_),
    .Y(_01745_));
 sky130_fd_sc_hs__nand2_1 _07173_ (.A(net2966),
    .B(net3143),
    .Y(_01746_));
 sky130_fd_sc_hs__xnor2_1 _07174_ (.A(net3225),
    .B(_01746_),
    .Y(_01747_));
 sky130_fd_sc_hs__and2_1 _07175_ (.A(net2141),
    .B(net2147),
    .X(_01748_));
 sky130_fd_sc_hs__nand4_2 _07176_ (.A(_01743_),
    .B(_01745_),
    .C(_01747_),
    .D(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hs__nand3_1 _07177_ (.A(_01716_),
    .B(_01718_),
    .C(net2166),
    .Y(_01750_));
 sky130_fd_sc_hs__nor2_1 _07178_ (.A(_01744_),
    .B(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hs__nor2_1 _07179_ (.A(net2131),
    .B(_01751_),
    .Y(_01752_));
 sky130_fd_sc_hs__nand2_1 _07180_ (.A(_01742_),
    .B(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hs__o21ai_1 _07181_ (.A1(_01741_),
    .A2(_01751_),
    .B1(net2131),
    .Y(_01754_));
 sky130_fd_sc_hs__nand2_1 _07182_ (.A(_01753_),
    .B(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hs__nand3_1 _07183_ (.A(net2141),
    .B(net2147),
    .C(_01720_),
    .Y(_01756_));
 sky130_fd_sc_hs__xnor2_1 _07184_ (.A(net2889),
    .B(net2166),
    .Y(_01757_));
 sky130_fd_sc_hs__nand2_1 _07185_ (.A(net3799),
    .B(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hs__o21a_1 _07186_ (.A1(net2166),
    .A2(net3799),
    .B1(_01758_),
    .X(_01759_));
 sky130_fd_sc_hs__xnor2_1 _07187_ (.A(_01756_),
    .B(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hs__nand2_1 _07188_ (.A(_01760_),
    .B(_01742_),
    .Y(_01761_));
 sky130_fd_sc_hs__nand3_1 _07189_ (.A(_01740_),
    .B(_01759_),
    .C(_01741_),
    .Y(_01762_));
 sky130_fd_sc_hs__nand2_2 _07190_ (.A(_01761_),
    .B(_01762_),
    .Y(_01763_));
 sky130_fd_sc_hs__nor2_2 _07191_ (.A(_01763_),
    .B(_01755_),
    .Y(_01764_));
 sky130_fd_sc_hs__nand2_2 _07192_ (.A(_01764_),
    .B(_01749_),
    .Y(_01765_));
 sky130_fd_sc_hs__nand2_1 _07193_ (.A(_01753_),
    .B(net2130),
    .Y(_01766_));
 sky130_fd_sc_hs__nand2_2 _07194_ (.A(_01766_),
    .B(net2120),
    .Y(_01767_));
 sky130_fd_sc_hs__nand2_2 _07195_ (.A(_01767_),
    .B(_01765_),
    .Y(_01768_));
 sky130_fd_sc_hs__nand2_2 _07196_ (.A(_01768_),
    .B(_01747_),
    .Y(_01769_));
 sky130_fd_sc_hs__inv_1 _07197_ (.A(_01747_),
    .Y(_01770_));
 sky130_fd_sc_hs__nand3_1 _07198_ (.A(_01765_),
    .B(_01770_),
    .C(_01767_),
    .Y(_01771_));
 sky130_fd_sc_hs__inv_1 _07199_ (.A(net3229),
    .Y(_01772_));
 sky130_fd_sc_hs__a21oi_1 _07200_ (.A1(net3230),
    .A2(net3180),
    .B1(net2945),
    .Y(_01773_));
 sky130_fd_sc_hs__xnor2_1 _07201_ (.A(_01772_),
    .B(_01773_),
    .Y(_01774_));
 sky130_fd_sc_hs__and2_2 _07202_ (.A(net3805),
    .B(_01745_),
    .X(_01775_));
 sky130_fd_sc_hs__nand4_4 _07203_ (.A(_01769_),
    .B(_01771_),
    .C(_01774_),
    .D(net2090),
    .Y(_01776_));
 sky130_fd_sc_hs__nand2_1 _07204_ (.A(_01775_),
    .B(_01747_),
    .Y(_01777_));
 sky130_fd_sc_hs__inv_1 _07205_ (.A(_01748_),
    .Y(_01778_));
 sky130_fd_sc_hs__nand2_1 _07206_ (.A(net3797),
    .B(_01778_),
    .Y(_01779_));
 sky130_fd_sc_hs__nand3_1 _07207_ (.A(net2114),
    .B(_01720_),
    .C(_01748_),
    .Y(_01780_));
 sky130_fd_sc_hs__and2_2 _07208_ (.A(_01779_),
    .B(_01780_),
    .X(_01781_));
 sky130_fd_sc_hs__nand2_1 _07209_ (.A(_01781_),
    .B(_01777_),
    .Y(_01782_));
 sky130_fd_sc_hs__nand4_1 _07210_ (.A(net2105),
    .B(net2112),
    .C(_01747_),
    .D(net2123),
    .Y(_01783_));
 sky130_fd_sc_hs__nand2_2 _07211_ (.A(_01782_),
    .B(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hs__nand2_1 _07212_ (.A(_01768_),
    .B(_01784_),
    .Y(_01785_));
 sky130_fd_sc_hs__nand3_1 _07213_ (.A(_01765_),
    .B(_01767_),
    .C(_01781_),
    .Y(_01786_));
 sky130_fd_sc_hs__nand2_2 _07214_ (.A(_01785_),
    .B(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hs__nand3_1 _07215_ (.A(_01743_),
    .B(net2113),
    .C(_01748_),
    .Y(_01788_));
 sky130_fd_sc_hs__nor2_1 _07216_ (.A(_01770_),
    .B(_01788_),
    .Y(_01789_));
 sky130_fd_sc_hs__nand2_1 _07217_ (.A(_01789_),
    .B(net2092),
    .Y(_01790_));
 sky130_fd_sc_hs__inv_1 _07218_ (.A(_01763_),
    .Y(_01791_));
 sky130_fd_sc_hs__nand2_1 _07219_ (.A(_01749_),
    .B(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hs__nand2_1 _07220_ (.A(_01790_),
    .B(net2086),
    .Y(_01793_));
 sky130_fd_sc_hs__nand2_2 _07221_ (.A(_01793_),
    .B(_01768_),
    .Y(_01794_));
 sky130_fd_sc_hs__nand2_1 _07222_ (.A(_01767_),
    .B(net2092),
    .Y(_01795_));
 sky130_fd_sc_hs__nand2_2 _07223_ (.A(_01794_),
    .B(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hs__nor2_4 _07224_ (.A(_01796_),
    .B(_01787_),
    .Y(_01797_));
 sky130_fd_sc_hs__nand2_2 _07225_ (.A(_01797_),
    .B(_01776_),
    .Y(_01798_));
 sky130_fd_sc_hs__o21ai_1 _07226_ (.A1(_01767_),
    .A2(_01792_),
    .B1(net2093),
    .Y(_01799_));
 sky130_fd_sc_hs__and2_1 _07227_ (.A(_01799_),
    .B(net4892),
    .X(_01800_));
 sky130_fd_sc_hs__inv_1 _07228_ (.A(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hs__nand3_2 _07229_ (.A(_01798_),
    .B(_01774_),
    .C(net2056),
    .Y(_01802_));
 sky130_fd_sc_hs__inv_1 _07230_ (.A(_01774_),
    .Y(_01803_));
 sky130_fd_sc_hs__o21ai_2 _07231_ (.A1(net2067),
    .A2(_01797_),
    .B1(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hs__nand2_2 _07232_ (.A(_01802_),
    .B(_01804_),
    .Y(_01805_));
 sky130_fd_sc_hs__inv_1 _07233_ (.A(net3230),
    .Y(_01806_));
 sky130_fd_sc_hs__nor2_1 _07234_ (.A(net3189),
    .B(net2945),
    .Y(_01807_));
 sky130_fd_sc_hs__xnor2_1 _07235_ (.A(_01806_),
    .B(_01807_),
    .Y(_01808_));
 sky130_fd_sc_hs__nand2_1 _07236_ (.A(net2068),
    .B(net2074),
    .Y(_01809_));
 sky130_fd_sc_hs__clkdlyinv3sd1_1 _07237_ (.A(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hs__nand3_2 _07238_ (.A(_01810_),
    .B(_01808_),
    .C(_01805_),
    .Y(_01811_));
 sky130_fd_sc_hs__and2_1 _07239_ (.A(net2091),
    .B(net2120),
    .X(_01812_));
 sky130_fd_sc_hs__o21ai_1 _07240_ (.A1(_01812_),
    .A2(_01764_),
    .B1(net2094),
    .Y(_01813_));
 sky130_fd_sc_hs__nand2_1 _07241_ (.A(_01813_),
    .B(net2088),
    .Y(_01814_));
 sky130_fd_sc_hs__nand3_1 _07242_ (.A(net2094),
    .B(_01812_),
    .C(net2092),
    .Y(_01815_));
 sky130_fd_sc_hs__nand2_1 _07243_ (.A(_01814_),
    .B(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hs__clkinv_2 _07244_ (.A(_01787_),
    .Y(_01817_));
 sky130_fd_sc_hs__o211ai_1 _07245_ (.A1(_01816_),
    .A2(_01800_),
    .B1(_01817_),
    .C1(net2058),
    .Y(_01818_));
 sky130_fd_sc_hs__a21o_1 _07246_ (.A1(_01776_),
    .A2(_01800_),
    .B1(_01817_),
    .X(_01819_));
 sky130_fd_sc_hs__nand2_1 _07247_ (.A(_01818_),
    .B(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hs__nand2_2 _07248_ (.A(net2056),
    .B(_01798_),
    .Y(_01821_));
 sky130_fd_sc_hs__nor2_1 _07249_ (.A(net2090),
    .B(_01768_),
    .Y(_01822_));
 sky130_fd_sc_hs__nand2_1 _07250_ (.A(net3796),
    .B(_01745_),
    .Y(_01823_));
 sky130_fd_sc_hs__xnor2_1 _07251_ (.A(_01770_),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hs__and2_2 _07252_ (.A(_01768_),
    .B(_01824_),
    .X(_01825_));
 sky130_fd_sc_hs__nor2_2 _07253_ (.A(_01822_),
    .B(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hs__nand3_1 _07254_ (.A(_01769_),
    .B(net2074),
    .C(_01774_),
    .Y(_01827_));
 sky130_fd_sc_hs__xnor2_1 _07255_ (.A(_01826_),
    .B(_01827_),
    .Y(_01828_));
 sky130_fd_sc_hs__nand2_1 _07256_ (.A(_01821_),
    .B(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hs__nand3_1 _07257_ (.A(_01798_),
    .B(net2056),
    .C(net2055),
    .Y(_01830_));
 sky130_fd_sc_hs__nand2_2 _07258_ (.A(_01830_),
    .B(_01829_),
    .Y(_01831_));
 sky130_fd_sc_hs__nor2_4 _07259_ (.A(_01831_),
    .B(_01820_),
    .Y(_01832_));
 sky130_fd_sc_hs__nand2_2 _07260_ (.A(_01832_),
    .B(_01811_),
    .Y(_01833_));
 sky130_fd_sc_hs__nand2_1 _07261_ (.A(_01776_),
    .B(_01817_),
    .Y(_01834_));
 sky130_fd_sc_hs__o21ai_1 _07262_ (.A1(_01801_),
    .A2(_01834_),
    .B1(net2057),
    .Y(_01835_));
 sky130_fd_sc_hs__and2_1 _07263_ (.A(_01835_),
    .B(net4902),
    .X(_01836_));
 sky130_fd_sc_hs__clkinv_1 _07264_ (.A(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hs__nand2_2 _07265_ (.A(_01837_),
    .B(_01833_),
    .Y(_01838_));
 sky130_fd_sc_hs__nand2_2 _07266_ (.A(_01838_),
    .B(_01808_),
    .Y(_01839_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _07267_ (.A(_01808_),
    .Y(_01840_));
 sky130_fd_sc_hs__nand3_2 _07268_ (.A(_01833_),
    .B(_01840_),
    .C(_01837_),
    .Y(_01841_));
 sky130_fd_sc_hs__nand2_1 _07269_ (.A(net2966),
    .B(net3224),
    .Y(_01842_));
 sky130_fd_sc_hs__xnor2_1 _07270_ (.A(net3232),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _07271_ (.A(_01843_),
    .Y(_01844_));
 sky130_fd_sc_hs__nand4_4 _07272_ (.A(_01839_),
    .B(_01841_),
    .C(_01844_),
    .D(net2028),
    .Y(_01845_));
 sky130_fd_sc_hs__and2_2 _07273_ (.A(net2041),
    .B(net2048),
    .X(_01846_));
 sky130_fd_sc_hs__nor2_2 _07274_ (.A(_01840_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hs__xnor2_1 _07275_ (.A(_01803_),
    .B(_01809_),
    .Y(_01848_));
 sky130_fd_sc_hs__nand2_1 _07276_ (.A(net2038),
    .B(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hs__o21ai_1 _07277_ (.A1(net2051),
    .A2(net2039),
    .B1(_01849_),
    .Y(_01850_));
 sky130_fd_sc_hs__nand2_1 _07278_ (.A(_01847_),
    .B(_01850_),
    .Y(_01851_));
 sky130_fd_sc_hs__o21a_1 _07279_ (.A1(_01810_),
    .A2(_01821_),
    .B1(_01849_),
    .X(_01852_));
 sky130_fd_sc_hs__nand2_1 _07280_ (.A(net2028),
    .B(_01808_),
    .Y(_01853_));
 sky130_fd_sc_hs__nand2_1 _07281_ (.A(_01852_),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hs__nand2_1 _07282_ (.A(_01851_),
    .B(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hs__nand2_1 _07283_ (.A(_01838_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hs__nand3_1 _07284_ (.A(_01833_),
    .B(_01852_),
    .C(_01837_),
    .Y(_01857_));
 sky130_fd_sc_hs__nand2_1 _07285_ (.A(_01856_),
    .B(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hs__inv_1 _07286_ (.A(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hs__inv_1 _07287_ (.A(net2014),
    .Y(_01860_));
 sky130_fd_sc_hs__nand2_1 _07288_ (.A(net2015),
    .B(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hs__nand2_1 _07289_ (.A(_01861_),
    .B(net2040),
    .Y(_01862_));
 sky130_fd_sc_hs__nand3_1 _07290_ (.A(_01862_),
    .B(net2027),
    .C(_01833_),
    .Y(_01863_));
 sky130_fd_sc_hs__and2_1 _07291_ (.A(_01818_),
    .B(_01819_),
    .X(_01864_));
 sky130_fd_sc_hs__nand3_1 _07292_ (.A(_01861_),
    .B(net2013),
    .C(net2037),
    .Y(_01865_));
 sky130_fd_sc_hs__nand2_2 _07293_ (.A(_01865_),
    .B(_01863_),
    .Y(_01866_));
 sky130_fd_sc_hs__o21ai_1 _07294_ (.A1(net2026),
    .A2(_01832_),
    .B1(_01811_),
    .Y(_01867_));
 sky130_fd_sc_hs__nand2_1 _07295_ (.A(_01867_),
    .B(net2014),
    .Y(_01868_));
 sky130_fd_sc_hs__o211ai_1 _07296_ (.A1(_01864_),
    .A2(net2026),
    .B1(_01860_),
    .C1(net2015),
    .Y(_01869_));
 sky130_fd_sc_hs__nand2_1 _07297_ (.A(_01868_),
    .B(_01869_),
    .Y(_01870_));
 sky130_fd_sc_hs__nand4_1 _07298_ (.A(net1971),
    .B(_01859_),
    .C(net1970),
    .D(net1983),
    .Y(_01871_));
 sky130_fd_sc_hs__nand2_1 _07299_ (.A(net1972),
    .B(_01859_),
    .Y(_01872_));
 sky130_fd_sc_hs__and2_1 _07300_ (.A(_01868_),
    .B(_01869_),
    .X(_01873_));
 sky130_fd_sc_hs__nand2_1 _07301_ (.A(_01872_),
    .B(net1982),
    .Y(_01874_));
 sky130_fd_sc_hs__nand2_2 _07302_ (.A(_01871_),
    .B(_01874_),
    .Y(_01875_));
 sky130_fd_sc_hs__o211ai_1 _07303_ (.A1(_01873_),
    .A2(net1969),
    .B1(_01859_),
    .C1(net1972),
    .Y(_01876_));
 sky130_fd_sc_hs__a21o_1 _07304_ (.A1(net1971),
    .A2(net4931),
    .B1(_01859_),
    .X(_01877_));
 sky130_fd_sc_hs__nand2_2 _07305_ (.A(_01877_),
    .B(_01876_),
    .Y(_01878_));
 sky130_fd_sc_hs__nor2_2 _07306_ (.A(_01870_),
    .B(_01858_),
    .Y(_01879_));
 sky130_fd_sc_hs__nand2_2 _07307_ (.A(_01879_),
    .B(_01845_),
    .Y(_01880_));
 sky130_fd_sc_hs__inv_2 _07308_ (.A(_01866_),
    .Y(_01881_));
 sky130_fd_sc_hs__nand2_2 _07309_ (.A(_01880_),
    .B(_01881_),
    .Y(_01882_));
 sky130_fd_sc_hs__nand2_1 _07310_ (.A(_01839_),
    .B(net2025),
    .Y(_01883_));
 sky130_fd_sc_hs__nand2_1 _07311_ (.A(net1991),
    .B(net2012),
    .Y(_01884_));
 sky130_fd_sc_hs__and2_2 _07312_ (.A(_01883_),
    .B(_01884_),
    .X(_01885_));
 sky130_fd_sc_hs__nand3_1 _07313_ (.A(net3835),
    .B(_01841_),
    .C(_01844_),
    .Y(_01886_));
 sky130_fd_sc_hs__nand2_1 _07314_ (.A(_01885_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hs__nand4_1 _07315_ (.A(net3834),
    .B(net1990),
    .C(_01844_),
    .D(net2025),
    .Y(_01888_));
 sky130_fd_sc_hs__nand2_2 _07316_ (.A(_01887_),
    .B(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hs__nand2_2 _07317_ (.A(_01882_),
    .B(_01889_),
    .Y(_01890_));
 sky130_fd_sc_hs__nand3_1 _07318_ (.A(_01880_),
    .B(_01885_),
    .C(_01881_),
    .Y(_01891_));
 sky130_fd_sc_hs__nand2_2 _07319_ (.A(_01890_),
    .B(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hs__nor2_4 _07320_ (.A(_01878_),
    .B(_01892_),
    .Y(_01893_));
 sky130_fd_sc_hs__nand2_2 _07321_ (.A(_01882_),
    .B(_01844_),
    .Y(_01894_));
 sky130_fd_sc_hs__nand3_2 _07322_ (.A(_01880_),
    .B(_01843_),
    .C(_01881_),
    .Y(_01895_));
 sky130_fd_sc_hs__nor2_1 _07323_ (.A(net3270),
    .B(net2945),
    .Y(_01896_));
 sky130_fd_sc_hs__xnor2_1 _07324_ (.A(net3308),
    .B(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _07325_ (.A(_01897_),
    .Y(_01898_));
 sky130_fd_sc_hs__nand2_2 _07326_ (.A(net3836),
    .B(_01841_),
    .Y(_01899_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _07327_ (.A(_01899_),
    .Y(_01900_));
 sky130_fd_sc_hs__nand4_2 _07328_ (.A(_01895_),
    .B(_01894_),
    .C(_01898_),
    .D(_01900_),
    .Y(_01901_));
 sky130_fd_sc_hs__o211ai_1 _07329_ (.A1(_01875_),
    .A2(_01893_),
    .B1(net1931),
    .C1(net3794),
    .Y(_01902_));
 sky130_fd_sc_hs__o21ai_1 _07330_ (.A1(net1942),
    .A2(_01893_),
    .B1(net3794),
    .Y(_01903_));
 sky130_fd_sc_hs__and2_1 _07331_ (.A(_01890_),
    .B(_01891_),
    .X(_01904_));
 sky130_fd_sc_hs__nand2_1 _07332_ (.A(_01903_),
    .B(net1929),
    .Y(_01905_));
 sky130_fd_sc_hs__nand2_2 _07333_ (.A(_01902_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hs__xnor2_1 _07334_ (.A(_01843_),
    .B(_01899_),
    .Y(_01907_));
 sky130_fd_sc_hs__nand2_1 _07335_ (.A(_01882_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hs__nand3_1 _07336_ (.A(net3803),
    .B(net1967),
    .C(_01881_),
    .Y(_01909_));
 sky130_fd_sc_hs__nand2_1 _07337_ (.A(_01908_),
    .B(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hs__nor2_1 _07338_ (.A(_01910_),
    .B(_01892_),
    .Y(_01911_));
 sky130_fd_sc_hs__nand2_2 _07339_ (.A(_01894_),
    .B(_01895_),
    .Y(_01912_));
 sky130_fd_sc_hs__nor2_1 _07340_ (.A(_01898_),
    .B(_01912_),
    .Y(_01913_));
 sky130_fd_sc_hs__nand2_1 _07341_ (.A(_01911_),
    .B(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hs__o21ai_1 _07342_ (.A1(net1968),
    .A2(_01912_),
    .B1(_01904_),
    .Y(_01915_));
 sky130_fd_sc_hs__nand2_1 _07343_ (.A(_01914_),
    .B(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hs__nand3_1 _07344_ (.A(_01916_),
    .B(net1950),
    .C(net1941),
    .Y(_01917_));
 sky130_fd_sc_hs__nand3b_1 _07345_ (.A_N(net1950),
    .B(_01914_),
    .C(_01915_),
    .Y(_01918_));
 sky130_fd_sc_hs__nand2_1 _07346_ (.A(_01917_),
    .B(_01918_),
    .Y(_01919_));
 sky130_fd_sc_hs__nor2_1 _07347_ (.A(_01906_),
    .B(_01919_),
    .Y(_01920_));
 sky130_fd_sc_hs__nand2_2 _07348_ (.A(_01901_),
    .B(_01893_),
    .Y(_01921_));
 sky130_fd_sc_hs__clkinv_1 _07349_ (.A(_01875_),
    .Y(_01922_));
 sky130_fd_sc_hs__nand2_2 _07350_ (.A(_01921_),
    .B(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hs__nand2_1 _07351_ (.A(net1927),
    .B(_01897_),
    .Y(_01924_));
 sky130_fd_sc_hs__nand3_1 _07352_ (.A(net1940),
    .B(net1949),
    .C(_01898_),
    .Y(_01925_));
 sky130_fd_sc_hs__nand2_1 _07353_ (.A(_01924_),
    .B(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hs__nand2_1 _07354_ (.A(_01923_),
    .B(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hs__nand3_1 _07355_ (.A(_01921_),
    .B(net1927),
    .C(_01922_),
    .Y(_01928_));
 sky130_fd_sc_hs__nand2_2 _07356_ (.A(_01927_),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hs__nand2_1 _07357_ (.A(_01925_),
    .B(net1928),
    .Y(_01930_));
 sky130_fd_sc_hs__nand2_1 _07358_ (.A(_01930_),
    .B(net1930),
    .Y(_01931_));
 sky130_fd_sc_hs__nand2_2 _07359_ (.A(_01923_),
    .B(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hs__nand3_1 _07360_ (.A(_01921_),
    .B(net1928),
    .C(_01922_),
    .Y(_01933_));
 sky130_fd_sc_hs__nand2_2 _07361_ (.A(_01933_),
    .B(_01932_),
    .Y(_01934_));
 sky130_fd_sc_hs__nor2_2 _07362_ (.A(_01929_),
    .B(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hs__nand2_1 _07363_ (.A(net2966),
    .B(net3390),
    .Y(_01936_));
 sky130_fd_sc_hs__xnor2_1 _07364_ (.A(net3307),
    .B(_01936_),
    .Y(_01937_));
 sky130_fd_sc_hs__nor2_1 _07365_ (.A(net3362),
    .B(net2945),
    .Y(_01938_));
 sky130_fd_sc_hs__xnor2_1 _07366_ (.A(net3459),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hs__nor2b_1 _07367_ (.A(_01939_),
    .B_N(_00154_),
    .Y(_01940_));
 sky130_fd_sc_hs__nand2_1 _07368_ (.A(_01940_),
    .B(net3672),
    .Y(_01941_));
 sky130_fd_sc_hs__or2_1 _07369_ (.A(_01937_),
    .B(_01941_),
    .X(_01942_));
 sky130_fd_sc_hs__nand2_2 _07370_ (.A(_01923_),
    .B(_01898_),
    .Y(_01943_));
 sky130_fd_sc_hs__nand3_1 _07371_ (.A(_01921_),
    .B(_01897_),
    .C(_01922_),
    .Y(_01944_));
 sky130_fd_sc_hs__nand2_2 _07372_ (.A(_01944_),
    .B(_01943_),
    .Y(_01945_));
 sky130_fd_sc_hs__nor2_2 _07373_ (.A(_01942_),
    .B(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hs__nand3_1 _07374_ (.A(_01920_),
    .B(_01935_),
    .C(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hs__buf_2 place2171 (.A(_05450_),
    .X(net2171));
 sky130_fd_sc_hs__nand2_2 _07376_ (.A(_01947_),
    .B(net2966),
    .Y(_01949_));
 sky130_fd_sc_hs__inv_1 _07377_ (.A(\u_window_buffer.write_ptr[27] ),
    .Y(_01950_));
 sky130_fd_sc_hs__nand2_1 _07378_ (.A(net1868),
    .B(net3670),
    .Y(_01951_));
 sky130_fd_sc_hs__buf_1 place2170 (.A(_05462_),
    .X(net2170));
 sky130_fd_sc_hs__buf_1 place2169 (.A(_05489_),
    .X(net2169));
 sky130_fd_sc_hs__nand3_1 _07381_ (.A(net1876),
    .B(net3691),
    .C(net2966),
    .Y(_01954_));
 sky130_fd_sc_hs__nand2_1 _07382_ (.A(_01951_),
    .B(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hs__nor2_4 _07383_ (.A(_01934_),
    .B(_01906_),
    .Y(_01956_));
 sky130_fd_sc_hs__nor2_1 _07384_ (.A(_01937_),
    .B(_01939_),
    .Y(_01957_));
 sky130_fd_sc_hs__nand2_1 _07385_ (.A(_01957_),
    .B(_00155_),
    .Y(_01958_));
 sky130_fd_sc_hs__or2_1 _07386_ (.A(_01958_),
    .B(net1927),
    .X(_01959_));
 sky130_fd_sc_hs__nor2_4 _07387_ (.A(_01945_),
    .B(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hs__and2_1 _07388_ (.A(_01917_),
    .B(_01918_),
    .X(_01961_));
 sky130_fd_sc_hs__nand3_2 _07389_ (.A(_01960_),
    .B(_01961_),
    .C(_01956_),
    .Y(_01962_));
 sky130_fd_sc_hs__nand2_8 _07390_ (.A(net3787),
    .B(net2966),
    .Y(_01963_));
 sky130_fd_sc_hs__buf_1 place2168 (.A(_01702_),
    .X(net2168));
 sky130_fd_sc_hs__inv_2 _07392_ (.A(\u_window_buffer.write_ptr[26] ),
    .Y(_01965_));
 sky130_fd_sc_hs__nand2_1 _07393_ (.A(_01963_),
    .B(net3668),
    .Y(_01966_));
 sky130_fd_sc_hs__buf_1 place2167 (.A(_01710_),
    .X(net2167));
 sky130_fd_sc_hs__buf_1 place2172 (.A(_05443_),
    .X(net2172));
 sky130_fd_sc_hs__nand3_1 _07396_ (.A(net1875),
    .B(net3692),
    .C(net2966),
    .Y(_01969_));
 sky130_fd_sc_hs__nand2_1 _07397_ (.A(_01966_),
    .B(_01969_),
    .Y(_01970_));
 sky130_fd_sc_hs__nand2_1 _07398_ (.A(_01955_),
    .B(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hs__nand2_1 _07399_ (.A(net1884),
    .B(_01946_),
    .Y(_01972_));
 sky130_fd_sc_hs__nand2_4 _07400_ (.A(_01972_),
    .B(net2966),
    .Y(_01973_));
 sky130_fd_sc_hs__o21ai_2 _07401_ (.A1(net1903),
    .A2(net1891),
    .B1(net2966),
    .Y(_01974_));
 sky130_fd_sc_hs__nand3_1 _07402_ (.A(_01973_),
    .B(net3693),
    .C(net1880),
    .Y(_01975_));
 sky130_fd_sc_hs__inv_1 _07403_ (.A(\u_window_buffer.write_ptr[25] ),
    .Y(_01976_));
 sky130_fd_sc_hs__nand3_1 _07404_ (.A(net1876),
    .B(net3666),
    .C(net2966),
    .Y(_01977_));
 sky130_fd_sc_hs__and2_1 _07405_ (.A(_01975_),
    .B(_01977_),
    .X(_01978_));
 sky130_fd_sc_hs__nand2_1 _07406_ (.A(net4934),
    .B(net3694),
    .Y(_01979_));
 sky130_fd_sc_hs__inv_1 _07407_ (.A(\u_window_buffer.write_ptr[24] ),
    .Y(_01980_));
 sky130_fd_sc_hs__nand3_1 _07408_ (.A(net1875),
    .B(net3665),
    .C(net2966),
    .Y(_01981_));
 sky130_fd_sc_hs__and2_2 _07409_ (.A(_01979_),
    .B(_01981_),
    .X(_01982_));
 sky130_fd_sc_hs__nand2_1 _07410_ (.A(_01978_),
    .B(_01982_),
    .Y(_01983_));
 sky130_fd_sc_hs__nor2_1 _07411_ (.A(_01971_),
    .B(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hs__inv_1 _07412_ (.A(\u_window_buffer.write_ptr[31] ),
    .Y(_01985_));
 sky130_fd_sc_hs__nand3_1 _07413_ (.A(_01973_),
    .B(net3664),
    .C(_01974_),
    .Y(_01986_));
 sky130_fd_sc_hs__nand3_1 _07414_ (.A(net1876),
    .B(net3685),
    .C(net2966),
    .Y(_01987_));
 sky130_fd_sc_hs__nand2_1 _07415_ (.A(_01986_),
    .B(_01987_),
    .Y(_01988_));
 sky130_fd_sc_hs__inv_1 _07416_ (.A(\u_window_buffer.write_ptr[30] ),
    .Y(_01989_));
 sky130_fd_sc_hs__nand2_1 _07417_ (.A(_01963_),
    .B(net3663),
    .Y(_01990_));
 sky130_fd_sc_hs__nand3_1 _07418_ (.A(net1875),
    .B(net3686),
    .C(net2966),
    .Y(_01991_));
 sky130_fd_sc_hs__nand2_2 _07419_ (.A(_01991_),
    .B(_01990_),
    .Y(_01992_));
 sky130_fd_sc_hs__nand2_1 _07420_ (.A(_01988_),
    .B(_01992_),
    .Y(_01993_));
 sky130_fd_sc_hs__inv_1 _07421_ (.A(net3689),
    .Y(_01994_));
 sky130_fd_sc_hs__nand2_1 _07422_ (.A(net1869),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hs__nand3_1 _07423_ (.A(net1876),
    .B(net3689),
    .C(net2966),
    .Y(_01996_));
 sky130_fd_sc_hs__nand2_1 _07424_ (.A(_01995_),
    .B(_01996_),
    .Y(_01997_));
 sky130_fd_sc_hs__inv_1 _07425_ (.A(net3690),
    .Y(_01998_));
 sky130_fd_sc_hs__nand2_1 _07426_ (.A(_01963_),
    .B(_01998_),
    .Y(_01999_));
 sky130_fd_sc_hs__nand3_1 _07427_ (.A(net1875),
    .B(net3690),
    .C(net2966),
    .Y(_02000_));
 sky130_fd_sc_hs__nand2_2 _07428_ (.A(_02000_),
    .B(_01999_),
    .Y(_02001_));
 sky130_fd_sc_hs__nand2_1 _07429_ (.A(_01997_),
    .B(_02001_),
    .Y(_02002_));
 sky130_fd_sc_hs__nor2_1 _07430_ (.A(_01993_),
    .B(_02002_),
    .Y(_02003_));
 sky130_fd_sc_hs__nand2_1 _07431_ (.A(_01984_),
    .B(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hs__nand2_1 _07432_ (.A(net4934),
    .B(net3698),
    .Y(_02005_));
 sky130_fd_sc_hs__inv_1 _07433_ (.A(\u_window_buffer.write_ptr[22] ),
    .Y(_02006_));
 sky130_fd_sc_hs__nand3_1 _07434_ (.A(net1875),
    .B(net3662),
    .C(net2966),
    .Y(_02007_));
 sky130_fd_sc_hs__nand2_2 _07435_ (.A(_02005_),
    .B(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hs__nand2_1 _07436_ (.A(net1869),
    .B(net3696),
    .Y(_02009_));
 sky130_fd_sc_hs__inv_1 _07437_ (.A(net3696),
    .Y(_02010_));
 sky130_fd_sc_hs__nand3_1 _07438_ (.A(net1876),
    .B(_02010_),
    .C(net2966),
    .Y(_02011_));
 sky130_fd_sc_hs__nand2_1 _07439_ (.A(_02009_),
    .B(_02011_),
    .Y(_02012_));
 sky130_fd_sc_hs__nor2_1 _07440_ (.A(_02012_),
    .B(_02008_),
    .Y(_02013_));
 sky130_fd_sc_hs__nand2_2 _07441_ (.A(net1866),
    .B(net3701),
    .Y(_02014_));
 sky130_fd_sc_hs__inv_1 _07442_ (.A(\u_window_buffer.write_ptr[20] ),
    .Y(_02015_));
 sky130_fd_sc_hs__nand3_1 _07443_ (.A(net1875),
    .B(net3661),
    .C(net2966),
    .Y(_02016_));
 sky130_fd_sc_hs__nand2_2 _07444_ (.A(_02016_),
    .B(_02014_),
    .Y(_02017_));
 sky130_fd_sc_hs__nand2_1 _07445_ (.A(net1868),
    .B(net3700),
    .Y(_02018_));
 sky130_fd_sc_hs__inv_1 _07446_ (.A(\u_window_buffer.write_ptr[21] ),
    .Y(_02019_));
 sky130_fd_sc_hs__nand3_1 _07447_ (.A(net1876),
    .B(net3660),
    .C(net2966),
    .Y(_02020_));
 sky130_fd_sc_hs__nand2_1 _07448_ (.A(_02018_),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hs__nor2_4 _07449_ (.A(_02021_),
    .B(_02017_),
    .Y(_02022_));
 sky130_fd_sc_hs__and2_1 _07450_ (.A(_02013_),
    .B(_02022_),
    .X(_02023_));
 sky130_fd_sc_hs__nand3_1 _07451_ (.A(_01973_),
    .B(net3705),
    .C(net1881),
    .Y(_02024_));
 sky130_fd_sc_hs__inv_1 _07452_ (.A(\u_window_buffer.write_ptr[17] ),
    .Y(_02025_));
 sky130_fd_sc_hs__nand3_1 _07453_ (.A(net1876),
    .B(net3656),
    .C(net2966),
    .Y(_02026_));
 sky130_fd_sc_hs__and2_2 _07454_ (.A(_02024_),
    .B(_02026_),
    .X(_02027_));
 sky130_fd_sc_hs__inv_1 _07455_ (.A(\u_window_buffer.write_ptr[16] ),
    .Y(_02028_));
 sky130_fd_sc_hs__nand2_1 _07456_ (.A(net3786),
    .B(net3655),
    .Y(_02029_));
 sky130_fd_sc_hs__nand3_1 _07457_ (.A(net1875),
    .B(net3706),
    .C(net2966),
    .Y(_02030_));
 sky130_fd_sc_hs__nand2_1 _07458_ (.A(_02029_),
    .B(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hs__nand2_1 _07459_ (.A(_02027_),
    .B(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hs__nand3_1 _07460_ (.A(_01973_),
    .B(net3703),
    .C(_01974_),
    .Y(_02033_));
 sky130_fd_sc_hs__inv_1 _07461_ (.A(\u_window_buffer.write_ptr[19] ),
    .Y(_02034_));
 sky130_fd_sc_hs__nand3_1 _07462_ (.A(net1876),
    .B(net3654),
    .C(net2966),
    .Y(_02035_));
 sky130_fd_sc_hs__and2_1 _07463_ (.A(_02033_),
    .B(_02035_),
    .X(_02036_));
 sky130_fd_sc_hs__nand2_1 _07464_ (.A(net3786),
    .B(net3704),
    .Y(_02037_));
 sky130_fd_sc_hs__inv_1 _07465_ (.A(\u_window_buffer.write_ptr[18] ),
    .Y(_02038_));
 sky130_fd_sc_hs__nand3_1 _07466_ (.A(net1875),
    .B(net3651),
    .C(net2966),
    .Y(_02039_));
 sky130_fd_sc_hs__and2_2 _07467_ (.A(_02037_),
    .B(_02039_),
    .X(_02040_));
 sky130_fd_sc_hs__nand2_1 _07468_ (.A(_02036_),
    .B(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hs__nor2_1 _07469_ (.A(_02032_),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hs__nand2_1 _07470_ (.A(_02023_),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hs__nor2_2 _07471_ (.A(_02043_),
    .B(_02004_),
    .Y(_02044_));
 sky130_fd_sc_hs__nor2_1 _07472_ (.A(net2945),
    .B(net1882),
    .Y(_02045_));
 sky130_fd_sc_hs__xnor2_1 _07473_ (.A(net3681),
    .B(net1890),
    .Y(_02046_));
 sky130_fd_sc_hs__xnor2_1 _07474_ (.A(_02045_),
    .B(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hs__inv_2 _07475_ (.A(\u_window_buffer.write_ptr[7] ),
    .Y(_02048_));
 sky130_fd_sc_hs__xnor2_1 _07476_ (.A(net3649),
    .B(net1904),
    .Y(_02049_));
 sky130_fd_sc_hs__xnor2_1 _07477_ (.A(_02049_),
    .B(_01973_),
    .Y(_02050_));
 sky130_fd_sc_hs__nor2_1 _07478_ (.A(_02047_),
    .B(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hs__o21ai_1 _07479_ (.A1(_00156_),
    .A2(net2945),
    .B1(_00766_),
    .Y(_02052_));
 sky130_fd_sc_hs__xnor2_1 _07480_ (.A(net3713),
    .B(net3744),
    .Y(_02053_));
 sky130_fd_sc_hs__o21ai_1 _07481_ (.A1(net3702),
    .A2(_02052_),
    .B1(_02053_),
    .Y(_02054_));
 sky130_fd_sc_hs__nor2_1 _07482_ (.A(_00155_),
    .B(net2945),
    .Y(_02055_));
 sky130_fd_sc_hs__xnor2_1 _07483_ (.A(net3687),
    .B(_02055_),
    .Y(_02056_));
 sky130_fd_sc_hs__xnor2_1 _07484_ (.A(_02056_),
    .B(_01939_),
    .Y(_02057_));
 sky130_fd_sc_hs__inv_1 _07485_ (.A(\u_window_buffer.write_ptr[3] ),
    .Y(_02058_));
 sky130_fd_sc_hs__xnor2_1 _07486_ (.A(net3648),
    .B(_01937_),
    .Y(_02059_));
 sky130_fd_sc_hs__nand2_1 _07487_ (.A(_01941_),
    .B(net2966),
    .Y(_02060_));
 sky130_fd_sc_hs__xnor2_1 _07488_ (.A(_02059_),
    .B(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hs__a2111oi_1 _07489_ (.A1(net3702),
    .A2(_02052_),
    .B1(_02054_),
    .C1(_02057_),
    .D1(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hs__o21ai_1 _07490_ (.A1(_01942_),
    .A2(net1889),
    .B1(net2966),
    .Y(_02063_));
 sky130_fd_sc_hs__xnor2_1 _07491_ (.A(net3682),
    .B(_01929_),
    .Y(_02064_));
 sky130_fd_sc_hs__or2_1 _07492_ (.A(_02063_),
    .B(_02064_),
    .X(_02065_));
 sky130_fd_sc_hs__nand2_1 _07493_ (.A(_02064_),
    .B(_02063_),
    .Y(_02066_));
 sky130_fd_sc_hs__clkinv_1 _07494_ (.A(\u_window_buffer.write_ptr[4] ),
    .Y(_02067_));
 sky130_fd_sc_hs__nand2_1 _07495_ (.A(_01958_),
    .B(net2966),
    .Y(_02068_));
 sky130_fd_sc_hs__xnor2_1 _07496_ (.A(net3646),
    .B(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hs__xnor2_1 _07497_ (.A(_02069_),
    .B(net1889),
    .Y(_02070_));
 sky130_fd_sc_hs__a21oi_1 _07498_ (.A1(_02065_),
    .A2(_02066_),
    .B1(_02070_),
    .Y(_02071_));
 sky130_fd_sc_hs__nand3_1 _07499_ (.A(_02051_),
    .B(net2807),
    .C(_02071_),
    .Y(_02072_));
 sky130_fd_sc_hs__inv_1 _07500_ (.A(\u_window_buffer.write_ptr[15] ),
    .Y(_02073_));
 sky130_fd_sc_hs__nand2_1 _07501_ (.A(net1868),
    .B(net3645),
    .Y(_02074_));
 sky130_fd_sc_hs__nand3_1 _07502_ (.A(net1876),
    .B(net3707),
    .C(net2966),
    .Y(_02075_));
 sky130_fd_sc_hs__nand2_1 _07503_ (.A(_02074_),
    .B(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hs__inv_1 _07504_ (.A(\u_window_buffer.write_ptr[14] ),
    .Y(_02077_));
 sky130_fd_sc_hs__nand2_1 _07505_ (.A(_01963_),
    .B(net3644),
    .Y(_02078_));
 sky130_fd_sc_hs__nand3_1 _07506_ (.A(net1875),
    .B(net3708),
    .C(net2966),
    .Y(_02079_));
 sky130_fd_sc_hs__nand2_1 _07507_ (.A(_02078_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hs__nand2_1 _07508_ (.A(_02076_),
    .B(_02080_),
    .Y(_02081_));
 sky130_fd_sc_hs__nand2_2 _07509_ (.A(_01973_),
    .B(_01974_),
    .Y(_02082_));
 sky130_fd_sc_hs__nand2_1 _07510_ (.A(_02082_),
    .B(net3709),
    .Y(_02083_));
 sky130_fd_sc_hs__inv_2 _07511_ (.A(\u_window_buffer.write_ptr[13] ),
    .Y(_02084_));
 sky130_fd_sc_hs__nand2_1 _07512_ (.A(net1868),
    .B(net3641),
    .Y(_02085_));
 sky130_fd_sc_hs__nand2_1 _07513_ (.A(_02083_),
    .B(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hs__clkinv_1 _07514_ (.A(\u_window_buffer.write_ptr[12] ),
    .Y(_02087_));
 sky130_fd_sc_hs__nand2_1 _07515_ (.A(net1867),
    .B(net3639),
    .Y(_02088_));
 sky130_fd_sc_hs__nand3_1 _07516_ (.A(net1875),
    .B(net3710),
    .C(net2966),
    .Y(_02089_));
 sky130_fd_sc_hs__nand2_1 _07517_ (.A(_02088_),
    .B(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hs__nand2_1 _07518_ (.A(_02086_),
    .B(_02090_),
    .Y(_02091_));
 sky130_fd_sc_hs__nor2_2 _07519_ (.A(_02081_),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hs__nand2_1 _07520_ (.A(net1883),
    .B(net1882),
    .Y(_02093_));
 sky130_fd_sc_hs__nand2_1 _07521_ (.A(_02093_),
    .B(net2966),
    .Y(_02094_));
 sky130_fd_sc_hs__inv_1 _07522_ (.A(\u_window_buffer.write_ptr[8] ),
    .Y(_02095_));
 sky130_fd_sc_hs__nand2_1 _07523_ (.A(net1892),
    .B(net3638),
    .Y(_02096_));
 sky130_fd_sc_hs__nand3_1 _07524_ (.A(net1902),
    .B(net1914),
    .C(net3679),
    .Y(_02097_));
 sky130_fd_sc_hs__and2_1 _07525_ (.A(_02096_),
    .B(_02097_),
    .X(_02098_));
 sky130_fd_sc_hs__nand2_1 _07526_ (.A(_02094_),
    .B(_02098_),
    .Y(_02099_));
 sky130_fd_sc_hs__nand2_1 _07527_ (.A(_02096_),
    .B(_02097_),
    .Y(_02100_));
 sky130_fd_sc_hs__nand3_1 _07528_ (.A(_02100_),
    .B(_02093_),
    .C(net2966),
    .Y(_02101_));
 sky130_fd_sc_hs__nand2_2 _07529_ (.A(_02099_),
    .B(_02101_),
    .Y(_02102_));
 sky130_fd_sc_hs__nand2_1 _07530_ (.A(net1868),
    .B(net3676),
    .Y(_02103_));
 sky130_fd_sc_hs__inv_1 _07531_ (.A(\u_window_buffer.write_ptr[9] ),
    .Y(_02104_));
 sky130_fd_sc_hs__nand3_1 _07532_ (.A(net1876),
    .B(net3637),
    .C(net2966),
    .Y(_02105_));
 sky130_fd_sc_hs__nand3_1 _07533_ (.A(_02102_),
    .B(_02103_),
    .C(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hs__nand2_1 _07534_ (.A(_02082_),
    .B(net3711),
    .Y(_02107_));
 sky130_fd_sc_hs__inv_2 _07535_ (.A(\u_window_buffer.write_ptr[11] ),
    .Y(_02108_));
 sky130_fd_sc_hs__nand2_1 _07536_ (.A(net1868),
    .B(net3634),
    .Y(_02109_));
 sky130_fd_sc_hs__nand2_1 _07537_ (.A(_02107_),
    .B(_02109_),
    .Y(_02110_));
 sky130_fd_sc_hs__inv_2 _07538_ (.A(\u_window_buffer.write_ptr[10] ),
    .Y(_02111_));
 sky130_fd_sc_hs__nand2_1 _07539_ (.A(_01963_),
    .B(net3632),
    .Y(_02112_));
 sky130_fd_sc_hs__nand3_1 _07540_ (.A(net1875),
    .B(net3712),
    .C(net2966),
    .Y(_02113_));
 sky130_fd_sc_hs__nand2_1 _07541_ (.A(_02113_),
    .B(_02112_),
    .Y(_02114_));
 sky130_fd_sc_hs__nand2_1 _07542_ (.A(_02110_),
    .B(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hs__nor2_1 _07543_ (.A(_02106_),
    .B(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hs__nand2_2 _07544_ (.A(_02116_),
    .B(_02092_),
    .Y(_02117_));
 sky130_fd_sc_hs__nor2_4 _07545_ (.A(_02117_),
    .B(_02072_),
    .Y(_02118_));
 sky130_fd_sc_hs__nand2_2 _07546_ (.A(_02044_),
    .B(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hs__nand3_2 _07547_ (.A(_02119_),
    .B(\u_window_buffer.next_state_is_valid_to_read ),
    .C(_00564_),
    .Y(_02120_));
 sky130_fd_sc_hs__nand2_2 _07548_ (.A(_02120_),
    .B(\u_hamming_window.hamming_state[2] ),
    .Y(_02121_));
 sky130_fd_sc_hs__buf_8 place2166 (.A(_01721_),
    .X(net2166));
 sky130_fd_sc_hs__nand2_2 _07550_ (.A(_02121_),
    .B(_00668_),
    .Y(_02123_));
 sky130_fd_sc_hs__a21oi_4 _07551_ (.A1(_00589_),
    .A2(_00565_),
    .B1(_02123_),
    .Y(_00022_));
 sky130_fd_sc_hs__and2_1 _07552_ (.A(hamming_done),
    .B(\u_fft.fft_state[0] ),
    .X(_02124_));
 sky130_fd_sc_hs__nand2_1 _07553_ (.A(_00037_),
    .B(_00040_),
    .Y(_02125_));
 sky130_fd_sc_hs__nand2_1 _07554_ (.A(_00049_),
    .B(_00052_),
    .Y(_02126_));
 sky130_fd_sc_hs__inv_1 _07555_ (.A(\u_fft.sched[45] ),
    .Y(_02127_));
 sky130_fd_sc_hs__nand2_1 _07556_ (.A(_00053_),
    .B(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hs__a21oi_1 _07557_ (.A1(_02128_),
    .A2(_00057_),
    .B1(_00056_),
    .Y(_02129_));
 sky130_fd_sc_hs__a21oi_1 _07558_ (.A1(_00049_),
    .A2(_00051_),
    .B1(_00048_),
    .Y(_02130_));
 sky130_fd_sc_hs__o21ai_1 _07559_ (.A1(_02126_),
    .A2(_02129_),
    .B1(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hs__a21o_1 _07560_ (.A1(_02131_),
    .A2(_00046_),
    .B1(_00045_),
    .X(_02132_));
 sky130_fd_sc_hs__a21oi_1 _07561_ (.A1(_02132_),
    .A2(_00043_),
    .B1(_00042_),
    .Y(_02133_));
 sky130_fd_sc_hs__a21oi_1 _07562_ (.A1(_00037_),
    .A2(_00039_),
    .B1(_00036_),
    .Y(_02134_));
 sky130_fd_sc_hs__o21ai_1 _07563_ (.A1(_02125_),
    .A2(_02133_),
    .B1(_02134_),
    .Y(_02135_));
 sky130_fd_sc_hs__or4_1 _07564_ (.A(\u_fft.sched[0] ),
    .B(\u_fft.sched[29] ),
    .C(_05778_),
    .D(_05786_),
    .X(_02136_));
 sky130_fd_sc_hs__nand4_1 _07565_ (.A(_02135_),
    .B(_00031_),
    .C(_00034_),
    .D(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hs__and2_1 _07566_ (.A(_00033_),
    .B(_00031_),
    .X(_02138_));
 sky130_fd_sc_hs__o21ai_1 _07567_ (.A1(_00030_),
    .A2(_02138_),
    .B1(_02136_),
    .Y(_02139_));
 sky130_fd_sc_hs__nand2_1 _07568_ (.A(_02137_),
    .B(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hs__nand2_1 _07569_ (.A(_00066_),
    .B(_00069_),
    .Y(_02141_));
 sky130_fd_sc_hs__nand2_1 _07570_ (.A(_00078_),
    .B(_00081_),
    .Y(_02142_));
 sky130_fd_sc_hs__inv_1 _07571_ (.A(_00183_),
    .Y(_02143_));
 sky130_fd_sc_hs__a21oi_1 _07572_ (.A1(_02143_),
    .A2(_00088_),
    .B1(_00087_),
    .Y(_02144_));
 sky130_fd_sc_hs__a21oi_1 _07573_ (.A1(_00078_),
    .A2(_00080_),
    .B1(_00077_),
    .Y(_02145_));
 sky130_fd_sc_hs__o21ai_1 _07574_ (.A1(_02142_),
    .A2(_02144_),
    .B1(_02145_),
    .Y(_02146_));
 sky130_fd_sc_hs__a21o_1 _07575_ (.A1(_02146_),
    .A2(_00075_),
    .B1(_00074_),
    .X(_02147_));
 sky130_fd_sc_hs__a21oi_1 _07576_ (.A1(_02147_),
    .A2(_00072_),
    .B1(_00071_),
    .Y(_02148_));
 sky130_fd_sc_hs__a21oi_1 _07577_ (.A1(_00066_),
    .A2(_00068_),
    .B1(_00065_),
    .Y(_02149_));
 sky130_fd_sc_hs__o21ai_1 _07578_ (.A1(_02141_),
    .A2(_02148_),
    .B1(_02149_),
    .Y(_02150_));
 sky130_fd_sc_hs__nand2_1 _07579_ (.A(_05800_),
    .B(_05794_),
    .Y(_02151_));
 sky130_fd_sc_hs__nand2_1 _07580_ (.A(_02151_),
    .B(\u_fft.sched[39] ),
    .Y(_02152_));
 sky130_fd_sc_hs__nand4_1 _07581_ (.A(_02150_),
    .B(_00060_),
    .C(_00063_),
    .D(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hs__and2_1 _07582_ (.A(_00062_),
    .B(_00060_),
    .X(_02154_));
 sky130_fd_sc_hs__o21ai_1 _07583_ (.A1(_00059_),
    .A2(_02154_),
    .B1(_02152_),
    .Y(_02155_));
 sky130_fd_sc_hs__nand2_1 _07584_ (.A(_02153_),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hs__and2_1 _07585_ (.A(_02140_),
    .B(_02156_),
    .X(_02157_));
 sky130_fd_sc_hs__inv_1 _07586_ (.A(\u_fft.sched[44] ),
    .Y(_02158_));
 sky130_fd_sc_hs__inv_2 _07587_ (.A(\u_fft.sched[42] ),
    .Y(_00176_));
 sky130_fd_sc_hs__inv_1 _07588_ (.A(\u_fft.sched[41] ),
    .Y(_00170_));
 sky130_fd_sc_hs__inv_2 _07589_ (.A(\u_fft.sched[40] ),
    .Y(_00169_));
 sky130_fd_sc_hs__nor2_1 _07590_ (.A(\u_fft.sched[44] ),
    .B(\u_fft.sched[43] ),
    .Y(_02159_));
 sky130_fd_sc_hs__a41oi_1 _07591_ (.A1(_02158_),
    .A2(_00176_),
    .A3(_00170_),
    .A4(_00169_),
    .B1(_02159_),
    .Y(_02160_));
 sky130_fd_sc_hs__inv_2 _07592_ (.A(\u_fft.fft_state[2] ),
    .Y(_02161_));
 sky130_fd_sc_hs__a21oi_1 _07593_ (.A1(_02157_),
    .A2(_02160_),
    .B1(_02161_),
    .Y(_02162_));
 sky130_fd_sc_hs__o21a_1 _07594_ (.A1(_02124_),
    .A2(_02162_),
    .B1(net211),
    .X(_00011_));
 sky130_fd_sc_hs__inv_1 _07595_ (.A(\u_fft.fft_state[0] ),
    .Y(_02163_));
 sky130_fd_sc_hs__nor2_1 _07596_ (.A(hamming_done),
    .B(_02163_),
    .Y(_02164_));
 sky130_fd_sc_hs__inv_2 _07597_ (.A(\u_fft.fft_state[3] ),
    .Y(_02165_));
 sky130_fd_sc_hs__nand3b_1 _07598_ (.A_N(_02164_),
    .B(net211),
    .C(_02165_),
    .Y(_00009_));
 sky130_fd_sc_hs__nand2_1 _07599_ (.A(_02160_),
    .B(\u_fft.fft_state[2] ),
    .Y(_02166_));
 sky130_fd_sc_hs__inv_2 _07600_ (.A(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hs__nand2_1 _07601_ (.A(_02157_),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hs__nand2b_1 _07602_ (.A_N(\u_fft.power_ptr_stage4[9] ),
    .B(\fft_ptr[8] ),
    .Y(_02169_));
 sky130_fd_sc_hs__nor3_1 _07603_ (.A(\fft_ptr[7] ),
    .B(\fft_ptr[6] ),
    .C(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hs__nor2_1 _07604_ (.A(\fft_ptr[1] ),
    .B(\fft_ptr[0] ),
    .Y(_02171_));
 sky130_fd_sc_hs__nor2_1 _07605_ (.A(\fft_ptr[3] ),
    .B(\fft_ptr[2] ),
    .Y(_02172_));
 sky130_fd_sc_hs__nor2_1 _07606_ (.A(\fft_ptr[5] ),
    .B(\fft_ptr[4] ),
    .Y(_02173_));
 sky130_fd_sc_hs__nand4_1 _07607_ (.A(_02170_),
    .B(_02171_),
    .C(_02172_),
    .D(_02173_),
    .Y(_02174_));
 sky130_fd_sc_hs__nand2_1 _07608_ (.A(_02174_),
    .B(\u_fft.fft_state[1] ),
    .Y(_02175_));
 sky130_fd_sc_hs__buf_1 place2164 (.A(_03436_),
    .X(net2164));
 sky130_fd_sc_hs__a21oi_1 _07610_ (.A1(_02168_),
    .A2(net3338),
    .B1(net3780),
    .Y(_00010_));
 sky130_fd_sc_hs__a21o_1 _07611_ (.A1(start_move_auto),
    .A2(net209),
    .B1(net212),
    .X(_00000_));
 sky130_fd_sc_hs__nor3_1 _07612_ (.A(idle),
    .B(\u_window_buffer.current_state[3] ),
    .C(\u_window_buffer.current_state[2] ),
    .Y(_02177_));
 sky130_fd_sc_hs__inv_1 _07613_ (.A(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hs__nor3_1 _07614_ (.A(\u_window_buffer.current_state[0] ),
    .B(\u_window_buffer.current_state[4] ),
    .C(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hs__o21ai_1 _07615_ (.A1(_00664_),
    .A2(_02179_),
    .B1(_00556_),
    .Y(_02180_));
 sky130_fd_sc_hs__inv_2 _07616_ (.A(_00557_),
    .Y(_02181_));
 sky130_fd_sc_hs__a21oi_1 _07617_ (.A1(_00593_),
    .A2(_02181_),
    .B1(_00592_),
    .Y(_02182_));
 sky130_fd_sc_hs__nand2_1 _07618_ (.A(_02179_),
    .B(_02181_),
    .Y(_02183_));
 sky130_fd_sc_hs__o31ai_1 _07619_ (.A1(_02179_),
    .A2(_02182_),
    .A3(_00659_),
    .B1(_02183_),
    .Y(_02184_));
 sky130_fd_sc_hs__a21oi_1 _07620_ (.A1(_00660_),
    .A2(_02180_),
    .B1(_02184_),
    .Y(_02185_));
 sky130_fd_sc_hs__o22ai_1 _07621_ (.A1(_00613_),
    .A2(_00665_),
    .B1(net3316),
    .B2(_00657_),
    .Y(_02186_));
 sky130_fd_sc_hs__a31o_1 _07622_ (.A1(_02184_),
    .A2(_00660_),
    .A3(_02180_),
    .B1(_02186_),
    .X(_02187_));
 sky130_fd_sc_hs__o21a_1 _07623_ (.A1(_02185_),
    .A2(_02187_),
    .B1(net1848),
    .X(_00025_));
 sky130_fd_sc_hs__inv_1 _07624_ (.A(net3754),
    .Y(_00211_));
 sky130_fd_sc_hs__clkinv_8 _07625_ (.A(net3774),
    .Y(_02188_));
 sky130_fd_sc_hs__clkinv_2 _07626_ (.A(net3775),
    .Y(_02189_));
 sky130_fd_sc_hs__inv_2 _07627_ (.A(net3745),
    .Y(_02190_));
 sky130_fd_sc_hs__inv_2 _07628_ (.A(net3746),
    .Y(_02191_));
 sky130_fd_sc_hs__nor2_4 _07629_ (.A(_02190_),
    .B(_02191_),
    .Y(_02192_));
 sky130_fd_sc_hs__inv_2 _07630_ (.A(net3747),
    .Y(_02193_));
 sky130_fd_sc_hs__inv_2 _07631_ (.A(_00220_),
    .Y(_02194_));
 sky130_fd_sc_hs__nand2_2 _07632_ (.A(net3626),
    .B(_02194_),
    .Y(_02195_));
 sky130_fd_sc_hs__nand3_2 _07633_ (.A(_02195_),
    .B(_02192_),
    .C(net3776),
    .Y(_02196_));
 sky130_fd_sc_hs__nor3_4 _07634_ (.A(_02188_),
    .B(_02189_),
    .C(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hs__and2_1 _07635_ (.A(net3771),
    .B(net3773),
    .X(_02198_));
 sky130_fd_sc_hs__nand2_2 _07636_ (.A(net3301),
    .B(net3625),
    .Y(_02199_));
 sky130_fd_sc_hs__clkinv_1 _07637_ (.A(net3762),
    .Y(_02200_));
 sky130_fd_sc_hs__inv_2 _07638_ (.A(net3763),
    .Y(_02201_));
 sky130_fd_sc_hs__nor2_1 _07639_ (.A(_02200_),
    .B(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hs__inv_1 _07640_ (.A(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hs__clkinv_1 _07641_ (.A(net3764),
    .Y(_02204_));
 sky130_fd_sc_hs__clkinv_1 _07642_ (.A(net3766),
    .Y(_02205_));
 sky130_fd_sc_hs__nor2_1 _07643_ (.A(_02204_),
    .B(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hs__bufinv_8 _07644_ (.A(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hs__nor2_1 _07645_ (.A(net3388),
    .B(net3387),
    .Y(_02208_));
 sky130_fd_sc_hs__clkdlyinv3sd1_1 _07646_ (.A(net3767),
    .Y(_02209_));
 sky130_fd_sc_hs__bufinv_8 _07647_ (.A(net3768),
    .Y(_02210_));
 sky130_fd_sc_hs__nor2_1 _07648_ (.A(_02209_),
    .B(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hs__inv_1 _07649_ (.A(net3769),
    .Y(_02212_));
 sky130_fd_sc_hs__inv_1 _07650_ (.A(net3770),
    .Y(_02213_));
 sky130_fd_sc_hs__nor2_1 _07651_ (.A(_02212_),
    .B(_02213_),
    .Y(_02214_));
 sky130_fd_sc_hs__nand2_1 _07652_ (.A(net3446),
    .B(net3445),
    .Y(_02215_));
 sky130_fd_sc_hs__inv_2 _07653_ (.A(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hs__nand2_1 _07654_ (.A(_02208_),
    .B(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hs__clkdlyinv3sd1_1 _07655_ (.A(net3758),
    .Y(_02218_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _07656_ (.A(net3759),
    .Y(_02219_));
 sky130_fd_sc_hs__clkinv_1 _07657_ (.A(net3760),
    .Y(_02220_));
 sky130_fd_sc_hs__inv_1 _07658_ (.A(net3761),
    .Y(_02221_));
 sky130_fd_sc_hs__nor4_1 _07659_ (.A(_02218_),
    .B(_02219_),
    .C(_02220_),
    .D(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hs__clkinv_1 _07660_ (.A(net3756),
    .Y(_02223_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _07661_ (.A(net3757),
    .Y(_02224_));
 sky130_fd_sc_hs__nor2_1 _07662_ (.A(_02223_),
    .B(_02224_),
    .Y(_02225_));
 sky130_fd_sc_hs__nand4_1 _07663_ (.A(_02222_),
    .B(net3753),
    .C(net3755),
    .D(_02225_),
    .Y(_02226_));
 sky130_fd_sc_hs__nor3_1 _07664_ (.A(net3266),
    .B(_02217_),
    .C(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hs__or2_1 _07665_ (.A(net3752),
    .B(_02227_),
    .X(_02228_));
 sky130_fd_sc_hs__nand2_1 _07666_ (.A(_02227_),
    .B(net3752),
    .Y(_02229_));
 sky130_fd_sc_hs__nand2_4 _07667_ (.A(_02228_),
    .B(_02229_),
    .Y(_02230_));
 sky130_fd_sc_hs__buf_1 place2163 (.A(_03448_),
    .X(net2163));
 sky130_fd_sc_hs__inv_2 _07669_ (.A(_02230_),
    .Y(_02232_));
 sky130_fd_sc_hs__bufbuf_8 place2162 (.A(_03484_),
    .X(net2162));
 sky130_fd_sc_hs__buf_1 place2161 (.A(_04545_),
    .X(net2161));
 sky130_fd_sc_hs__nor2_1 _07672_ (.A(net3754),
    .B(net3090),
    .Y(_02235_));
 sky130_fd_sc_hs__o21bai_1 _07673_ (.A1(_00213_),
    .A2(net3132),
    .B1_N(_02235_),
    .Y(_00215_));
 sky130_fd_sc_hs__buf_1 place2160 (.A(_04555_),
    .X(net2160));
 sky130_fd_sc_hs__inv_1 _07675_ (.A(\u_hamming_window.hamming_state[1] ),
    .Y(_02237_));
 sky130_fd_sc_hs__nor3_1 _07676_ (.A(net3782),
    .B(_02237_),
    .C(_00588_),
    .Y(_00004_));
 sky130_fd_sc_hs__inv_1 _07677_ (.A(\u_dct.dct_state[2] ),
    .Y(_02238_));
 sky130_fd_sc_hs__nor3_1 _07678_ (.A(net3781),
    .B(_02238_),
    .C(_00571_),
    .Y(_00001_));
 sky130_fd_sc_hs__inv_1 _07679_ (.A(\u_dct.dct_state[1] ),
    .Y(_02239_));
 sky130_fd_sc_hs__nor3_1 _07680_ (.A(net3781),
    .B(_02239_),
    .C(_00573_),
    .Y(_00002_));
 sky130_fd_sc_hs__nor2_1 _07681_ (.A(_05815_),
    .B(_05822_),
    .Y(_00005_));
 sky130_fd_sc_hs__inv_1 _07682_ (.A(\u_fft.fft_state[1] ),
    .Y(_02240_));
 sky130_fd_sc_hs__nor3_1 _07683_ (.A(net3780),
    .B(_02240_),
    .C(_02174_),
    .Y(_00003_));
 sky130_fd_sc_hs__inv_1 _07684_ (.A(\u_dct.k_ptr[0] ),
    .Y(_00159_));
 sky130_fd_sc_hs__inv_1 _07685_ (.A(\u_dct.n_ptr[0] ),
    .Y(_00164_));
 sky130_fd_sc_hs__inv_2 _07686_ (.A(\mel_ptr[0] ),
    .Y(_00205_));
 sky130_fd_sc_hs__inv_2 _07687_ (.A(net3765),
    .Y(_00210_));
 sky130_fd_sc_hs__inv_1 _07688_ (.A(\u_window_buffer.move_counter[0] ),
    .Y(_00221_));
 sky130_fd_sc_hs__inv_1 _07689_ (.A(\u_hamming_window.calc_pointer[0] ),
    .Y(_00235_));
 sky130_fd_sc_hs__inv_2 _07690_ (.A(\u_mel.k[0] ),
    .Y(\u_mel.k_next[0] ));
 sky130_fd_sc_hs__inv_1 _07691_ (.A(\u_fft.sched[21] ),
    .Y(_00054_));
 sky130_fd_sc_hs__inv_1 _07692_ (.A(\u_dct.k_ptr[1] ),
    .Y(_00160_));
 sky130_fd_sc_hs__inv_1 _07693_ (.A(\u_dct.n_ptr[1] ),
    .Y(_00165_));
 sky130_fd_sc_hs__inv_2 _07694_ (.A(\u_fft.sched[55] ),
    .Y(_00182_));
 sky130_fd_sc_hs__inv_1 _07695_ (.A(\mel_ptr[1] ),
    .Y(_00206_));
 sky130_fd_sc_hs__inv_1 _07696_ (.A(\u_window_buffer.move_counter[1] ),
    .Y(_00222_));
 sky130_fd_sc_hs__inv_2 _07697_ (.A(\u_hamming_window.calc_pointer[1] ),
    .Y(_00236_));
 sky130_fd_sc_hs__inv_1 _07698_ (.A(\u_mel.k[1] ),
    .Y(_00240_));
 sky130_fd_sc_hs__inv_1 _07699_ (.A(_00085_),
    .Y(_00086_));
 sky130_fd_sc_hs__buf_1 place2158 (.A(_04569_),
    .X(net2158));
 sky130_fd_sc_hs__o21ai_1 _07701_ (.A1(hamming_done),
    .A2(hamming_finished),
    .B1(net3784),
    .Y(_02242_));
 sky130_fd_sc_hs__a21oi_1 _07702_ (.A1(hamming_finished),
    .A2(idle),
    .B1(_02242_),
    .Y(_00243_));
 sky130_fd_sc_hs__buf_1 place2165 (.A(_03436_),
    .X(net2165));
 sky130_fd_sc_hs__nor3b_1 _07704_ (.A(_05774_),
    .B(_00592_),
    .C_N(hamming_finished),
    .Y(_00244_));
 sky130_fd_sc_hs__nand2_1 _07705_ (.A(_00612_),
    .B(fifo_rd_en),
    .Y(_02244_));
 sky130_fd_sc_hs__o21ai_1 _07706_ (.A1(_00230_),
    .A2(_02244_),
    .B1(net211),
    .Y(_02245_));
 sky130_fd_sc_hs__a21oi_1 _07707_ (.A1(_00230_),
    .A2(_02244_),
    .B1(_02245_),
    .Y(_00245_));
 sky130_fd_sc_hs__o21ai_1 _07708_ (.A1(_00233_),
    .A2(_02244_),
    .B1(net211),
    .Y(_02246_));
 sky130_fd_sc_hs__a21oi_1 _07709_ (.A1(_00231_),
    .A2(_02244_),
    .B1(_02246_),
    .Y(_00246_));
 sky130_fd_sc_hs__inv_2 _07710_ (.A(_02244_),
    .Y(_02247_));
 sky130_fd_sc_hs__and2_1 _07711_ (.A(_02247_),
    .B(_00234_),
    .X(_02248_));
 sky130_fd_sc_hs__nor2_1 _07712_ (.A(\tx_fifo.read_ptr[2] ),
    .B(_02248_),
    .Y(_02249_));
 sky130_fd_sc_hs__nand2_1 _07713_ (.A(_02248_),
    .B(\tx_fifo.read_ptr[2] ),
    .Y(_02250_));
 sky130_fd_sc_hs__nor3b_1 _07714_ (.A(net3781),
    .B(_02249_),
    .C_N(_02250_),
    .Y(_00247_));
 sky130_fd_sc_hs__nor3_1 _07715_ (.A(_00230_),
    .B(_00231_),
    .C(_00598_),
    .Y(_02251_));
 sky130_fd_sc_hs__nor3b_1 _07716_ (.A(_00600_),
    .B(_02244_),
    .C_N(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hs__a21oi_1 _07717_ (.A1(_02247_),
    .A2(_02251_),
    .B1(\tx_fifo.read_ptr[3] ),
    .Y(_02253_));
 sky130_fd_sc_hs__nor3_1 _07718_ (.A(net3781),
    .B(_02252_),
    .C(_02253_),
    .Y(_00248_));
 sky130_fd_sc_hs__bufbuf_8 place2159 (.A(_04566_),
    .X(net2159));
 sky130_fd_sc_hs__nor2_1 _07720_ (.A(_00600_),
    .B(_02250_),
    .Y(_02255_));
 sky130_fd_sc_hs__nor2_1 _07721_ (.A(\tx_fifo.read_ptr[4] ),
    .B(_02255_),
    .Y(_02256_));
 sky130_fd_sc_hs__nand2_1 _07722_ (.A(_02255_),
    .B(\tx_fifo.read_ptr[4] ),
    .Y(_02257_));
 sky130_fd_sc_hs__nor3b_1 _07723_ (.A(net3781),
    .B(_02256_),
    .C_N(_02257_),
    .Y(_00249_));
 sky130_fd_sc_hs__clkinv_1 _07724_ (.A(\tx_fifo.read_ptr[5] ),
    .Y(_02258_));
 sky130_fd_sc_hs__nand2_1 _07725_ (.A(_02252_),
    .B(\tx_fifo.read_ptr[4] ),
    .Y(_02259_));
 sky130_fd_sc_hs__nor2_1 _07726_ (.A(_02258_),
    .B(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hs__inv_1 _07727_ (.A(_02260_),
    .Y(_02261_));
 sky130_fd_sc_hs__nand2_1 _07728_ (.A(_02261_),
    .B(net211),
    .Y(_02262_));
 sky130_fd_sc_hs__a21oi_1 _07729_ (.A1(_02258_),
    .A2(_02259_),
    .B1(_02262_),
    .Y(_00250_));
 sky130_fd_sc_hs__nor3_1 _07730_ (.A(_02258_),
    .B(_00603_),
    .C(_02257_),
    .Y(_02263_));
 sky130_fd_sc_hs__a31oi_1 _07731_ (.A1(_02255_),
    .A2(\tx_fifo.read_ptr[4] ),
    .A3(\tx_fifo.read_ptr[5] ),
    .B1(\tx_fifo.read_ptr[6] ),
    .Y(_02264_));
 sky130_fd_sc_hs__nor3_1 _07732_ (.A(net3781),
    .B(_02263_),
    .C(_02264_),
    .Y(_00251_));
 sky130_fd_sc_hs__a21oi_1 _07733_ (.A1(_02260_),
    .A2(\tx_fifo.read_ptr[6] ),
    .B1(\tx_fifo.read_ptr[7] ),
    .Y(_02265_));
 sky130_fd_sc_hs__inv_1 _07734_ (.A(\tx_fifo.read_ptr[7] ),
    .Y(_02266_));
 sky130_fd_sc_hs__nor3_1 _07735_ (.A(_00603_),
    .B(_02266_),
    .C(_02261_),
    .Y(_02267_));
 sky130_fd_sc_hs__nor3_1 _07736_ (.A(net3781),
    .B(_02265_),
    .C(_02267_),
    .Y(_00252_));
 sky130_fd_sc_hs__clkinv_1 _07737_ (.A(\tx_fifo.write_ptr[4] ),
    .Y(_02268_));
 sky130_fd_sc_hs__inv_1 _07738_ (.A(\tx_fifo.write_ptr[3] ),
    .Y(_02269_));
 sky130_fd_sc_hs__nand3_1 _07739_ (.A(\tx_fifo.write_ptr[0] ),
    .B(\tx_fifo.write_ptr[1] ),
    .C(\tx_fifo.write_ptr[2] ),
    .Y(_02270_));
 sky130_fd_sc_hs__nor2_1 _07740_ (.A(_02269_),
    .B(_02270_),
    .Y(_02271_));
 sky130_fd_sc_hs__inv_1 _07741_ (.A(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hs__nor2_1 _07742_ (.A(_02268_),
    .B(_02272_),
    .Y(_02273_));
 sky130_fd_sc_hs__inv_1 _07743_ (.A(\tx_fifo.write_ptr[5] ),
    .Y(_02274_));
 sky130_fd_sc_hs__nor2_1 _07744_ (.A(_02268_),
    .B(_02274_),
    .Y(_02275_));
 sky130_fd_sc_hs__inv_1 _07745_ (.A(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hs__inv_1 _07746_ (.A(\tx_fifo.write_ptr[2] ),
    .Y(_02277_));
 sky130_fd_sc_hs__inv_1 _07747_ (.A(_00157_),
    .Y(_02278_));
 sky130_fd_sc_hs__nor3_1 _07748_ (.A(_02277_),
    .B(_02269_),
    .C(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hs__inv_2 _07749_ (.A(_02279_),
    .Y(_02280_));
 sky130_fd_sc_hs__nor2_1 _07750_ (.A(_02276_),
    .B(_02280_),
    .Y(_02281_));
 sky130_fd_sc_hs__nand3_1 _07751_ (.A(_02275_),
    .B(\tx_fifo.write_ptr[6] ),
    .C(\tx_fifo.write_ptr[7] ),
    .Y(_02282_));
 sky130_fd_sc_hs__nor2_1 _07752_ (.A(_02282_),
    .B(_02280_),
    .Y(_02283_));
 sky130_fd_sc_hs__a21oi_1 _07753_ (.A1(_02281_),
    .A2(_00605_),
    .B1(_02283_),
    .Y(_02284_));
 sky130_fd_sc_hs__xnor2_1 _07754_ (.A(\tx_fifo.read_ptr[1] ),
    .B(_00158_),
    .Y(_02285_));
 sky130_fd_sc_hs__nand2_1 _07755_ (.A(_00609_),
    .B(_02285_),
    .Y(_02286_));
 sky130_fd_sc_hs__o22ai_1 _07756_ (.A1(_02278_),
    .A2(_00599_),
    .B1(_00595_),
    .B2(_02279_),
    .Y(_02287_));
 sky130_fd_sc_hs__nand2_1 _07757_ (.A(_00599_),
    .B(_02278_),
    .Y(_02288_));
 sky130_fd_sc_hs__nand2_1 _07758_ (.A(_02279_),
    .B(_00595_),
    .Y(_02289_));
 sky130_fd_sc_hs__o211ai_1 _07759_ (.A1(_02270_),
    .A2(_00601_),
    .B1(_02288_),
    .C1(_02289_),
    .Y(_02290_));
 sky130_fd_sc_hs__a2111oi_1 _07760_ (.A1(_00601_),
    .A2(_02270_),
    .B1(_02286_),
    .C1(_02287_),
    .D1(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hs__inv_1 _07761_ (.A(_02281_),
    .Y(_02292_));
 sky130_fd_sc_hs__inv_1 _07762_ (.A(\tx_fifo.write_ptr[6] ),
    .Y(_02293_));
 sky130_fd_sc_hs__nor4_1 _07763_ (.A(_02268_),
    .B(_02274_),
    .C(_02293_),
    .D(_02272_),
    .Y(_02294_));
 sky130_fd_sc_hs__xnor2_1 _07764_ (.A(_00606_),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hs__a221oi_1 _07765_ (.A1(_00604_),
    .A2(_02292_),
    .B1(_00596_),
    .B2(_02273_),
    .C1(_02295_),
    .Y(_02296_));
 sky130_fd_sc_hs__o2111ai_1 _07766_ (.A1(_00596_),
    .A2(_02273_),
    .B1(_02284_),
    .C1(_02291_),
    .D1(_02296_),
    .Y(_02297_));
 sky130_fd_sc_hs__nand3_1 _07767_ (.A(_00603_),
    .B(_02266_),
    .C(_00232_),
    .Y(_02298_));
 sky130_fd_sc_hs__or4_1 _07768_ (.A(\tx_fifo.read_ptr[2] ),
    .B(\tx_fifo.read_ptr[3] ),
    .C(\tx_fifo.read_ptr[4] ),
    .D(\tx_fifo.read_ptr[5] ),
    .X(_02299_));
 sky130_fd_sc_hs__o41a_1 _07769_ (.A1(_02280_),
    .A2(_02282_),
    .A3(_02298_),
    .A4(_02299_),
    .B1(pre_emphasis_valid),
    .X(_02300_));
 sky130_fd_sc_hs__nand2_1 _07770_ (.A(_02297_),
    .B(_02300_),
    .Y(_02301_));
 sky130_fd_sc_hs__inv_2 _07771_ (.A(_02301_),
    .Y(_02302_));
 sky130_fd_sc_hs__o21ai_1 _07772_ (.A1(\tx_fifo.write_ptr[0] ),
    .A2(_02302_),
    .B1(net211),
    .Y(_02303_));
 sky130_fd_sc_hs__a21oi_1 _07773_ (.A1(\tx_fifo.write_ptr[0] ),
    .A2(_02302_),
    .B1(_02303_),
    .Y(_00253_));
 sky130_fd_sc_hs__nand2_1 _07774_ (.A(_02302_),
    .B(_00158_),
    .Y(_02304_));
 sky130_fd_sc_hs__nand2_1 _07775_ (.A(_02301_),
    .B(\tx_fifo.write_ptr[1] ),
    .Y(_02305_));
 sky130_fd_sc_hs__a21oi_1 _07776_ (.A1(_02304_),
    .A2(_02305_),
    .B1(net3781),
    .Y(_00254_));
 sky130_fd_sc_hs__nor3_1 _07777_ (.A(_02277_),
    .B(_02278_),
    .C(_02301_),
    .Y(_02306_));
 sky130_fd_sc_hs__a21oi_1 _07778_ (.A1(_02302_),
    .A2(_00157_),
    .B1(\tx_fifo.write_ptr[2] ),
    .Y(_02307_));
 sky130_fd_sc_hs__nor3_1 _07779_ (.A(net3781),
    .B(_02306_),
    .C(_02307_),
    .Y(_00255_));
 sky130_fd_sc_hs__nor2_1 _07780_ (.A(_02272_),
    .B(_02301_),
    .Y(_02308_));
 sky130_fd_sc_hs__o21a_1 _07781_ (.A1(_02270_),
    .A2(_02301_),
    .B1(_02269_),
    .X(_02309_));
 sky130_fd_sc_hs__nor3_1 _07782_ (.A(net3781),
    .B(_02308_),
    .C(_02309_),
    .Y(_00256_));
 sky130_fd_sc_hs__nor3_1 _07783_ (.A(_02268_),
    .B(_02280_),
    .C(_02301_),
    .Y(_02310_));
 sky130_fd_sc_hs__a21oi_1 _07784_ (.A1(_02302_),
    .A2(_02279_),
    .B1(\tx_fifo.write_ptr[4] ),
    .Y(_02311_));
 sky130_fd_sc_hs__nor3_1 _07785_ (.A(net3781),
    .B(_02310_),
    .C(_02311_),
    .Y(_00257_));
 sky130_fd_sc_hs__a21oi_1 _07786_ (.A1(_02302_),
    .A2(_02273_),
    .B1(\tx_fifo.write_ptr[5] ),
    .Y(_02312_));
 sky130_fd_sc_hs__a211oi_1 _07787_ (.A1(_02275_),
    .A2(_02308_),
    .B1(net3781),
    .C1(_02312_),
    .Y(_00258_));
 sky130_fd_sc_hs__buf_1 place2156 (.A(_03465_),
    .X(net2156));
 sky130_fd_sc_hs__nor3_1 _07789_ (.A(_02293_),
    .B(_02292_),
    .C(_02301_),
    .Y(_02314_));
 sky130_fd_sc_hs__a21oi_1 _07790_ (.A1(_02302_),
    .A2(_02281_),
    .B1(\tx_fifo.write_ptr[6] ),
    .Y(_02315_));
 sky130_fd_sc_hs__nor3_1 _07791_ (.A(net3781),
    .B(_02314_),
    .C(_02315_),
    .Y(_00259_));
 sky130_fd_sc_hs__nor3_1 _07792_ (.A(_02282_),
    .B(_02272_),
    .C(_02301_),
    .Y(_02316_));
 sky130_fd_sc_hs__a21oi_1 _07793_ (.A1(_02302_),
    .A2(_02294_),
    .B1(\tx_fifo.write_ptr[7] ),
    .Y(_02317_));
 sky130_fd_sc_hs__nor3_1 _07794_ (.A(net3781),
    .B(_02316_),
    .C(_02317_),
    .Y(_00260_));
 sky130_fd_sc_hs__nor2_1 _07795_ (.A(net3781),
    .B(_00580_),
    .Y(_00261_));
 sky130_fd_sc_hs__a21oi_1 _07796_ (.A1(_02239_),
    .A2(_00577_),
    .B1(_00578_),
    .Y(_02318_));
 sky130_fd_sc_hs__nor2_1 _07797_ (.A(_02239_),
    .B(_00578_),
    .Y(_02319_));
 sky130_fd_sc_hs__nor2_1 _07798_ (.A(\u_dct.k_ptr[0] ),
    .B(_02319_),
    .Y(_02320_));
 sky130_fd_sc_hs__a211oi_1 _07799_ (.A1(net3386),
    .A2(\u_dct.k_ptr[0] ),
    .B1(net3781),
    .C1(_02320_),
    .Y(_00262_));
 sky130_fd_sc_hs__inv_2 _07800_ (.A(net3386),
    .Y(_02321_));
 sky130_fd_sc_hs__nand2_1 _07801_ (.A(_02321_),
    .B(\u_dct.k_ptr[1] ),
    .Y(_02322_));
 sky130_fd_sc_hs__nand2_1 _07802_ (.A(_02319_),
    .B(_00162_),
    .Y(_02323_));
 sky130_fd_sc_hs__buf_1 place2157 (.A(_03465_),
    .X(net2157));
 sky130_fd_sc_hs__a21oi_1 _07804_ (.A1(_02322_),
    .A2(_02323_),
    .B1(net3781),
    .Y(_00263_));
 sky130_fd_sc_hs__a21oi_1 _07805_ (.A1(net3386),
    .A2(_00163_),
    .B1(\u_dct.k_ptr[2] ),
    .Y(_02325_));
 sky130_fd_sc_hs__o21ai_1 _07806_ (.A1(\u_dct.dct_state[1] ),
    .A2(_00575_),
    .B1(net211),
    .Y(_02326_));
 sky130_fd_sc_hs__inv_1 _07807_ (.A(\u_dct.k_ptr[2] ),
    .Y(_02327_));
 sky130_fd_sc_hs__nor3b_1 _07808_ (.A(_02327_),
    .B(_02321_),
    .C_N(_00163_),
    .Y(_02328_));
 sky130_fd_sc_hs__nor3_1 _07809_ (.A(_02325_),
    .B(_02326_),
    .C(_02328_),
    .Y(_00264_));
 sky130_fd_sc_hs__nor3_1 _07810_ (.A(_02327_),
    .B(_00159_),
    .C(_00160_),
    .Y(_02329_));
 sky130_fd_sc_hs__and3_1 _07811_ (.A(net3386),
    .B(_02329_),
    .C(\u_dct.k_ptr[3] ),
    .X(_02330_));
 sky130_fd_sc_hs__a21oi_1 _07812_ (.A1(net3386),
    .A2(_02329_),
    .B1(\u_dct.k_ptr[3] ),
    .Y(_02331_));
 sky130_fd_sc_hs__nor3_1 _07813_ (.A(_02326_),
    .B(_02330_),
    .C(_02331_),
    .Y(_00265_));
 sky130_fd_sc_hs__nor2_1 _07814_ (.A(_02238_),
    .B(_00578_),
    .Y(_02332_));
 sky130_fd_sc_hs__nor2_1 _07815_ (.A(\u_dct.n_ptr[0] ),
    .B(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hs__nor2_1 _07816_ (.A(_02332_),
    .B(_02318_),
    .Y(_02334_));
 sky130_fd_sc_hs__nor2_1 _07817_ (.A(_00164_),
    .B(_02334_),
    .Y(_02335_));
 sky130_fd_sc_hs__nor3_1 _07818_ (.A(net3781),
    .B(_02333_),
    .C(_02335_),
    .Y(_00266_));
 sky130_fd_sc_hs__nand2_1 _07819_ (.A(_02334_),
    .B(\u_dct.n_ptr[1] ),
    .Y(_02336_));
 sky130_fd_sc_hs__nand2_1 _07820_ (.A(_02332_),
    .B(_00167_),
    .Y(_02337_));
 sky130_fd_sc_hs__a21oi_1 _07821_ (.A1(_02336_),
    .A2(_02337_),
    .B1(net3781),
    .Y(_00267_));
 sky130_fd_sc_hs__o21a_1 _07822_ (.A1(_02332_),
    .A2(net3386),
    .B1(_00168_),
    .X(_02338_));
 sky130_fd_sc_hs__nor2_1 _07823_ (.A(\u_dct.n_ptr[2] ),
    .B(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hs__o21ai_1 _07824_ (.A1(\u_dct.dct_state[2] ),
    .A2(_02321_),
    .B1(net211),
    .Y(_02340_));
 sky130_fd_sc_hs__nand2_1 _07825_ (.A(_02338_),
    .B(\u_dct.n_ptr[2] ),
    .Y(_02341_));
 sky130_fd_sc_hs__clkinv_1 _07826_ (.A(_02341_),
    .Y(_02342_));
 sky130_fd_sc_hs__nor3_1 _07827_ (.A(_02339_),
    .B(_02340_),
    .C(_02342_),
    .Y(_00268_));
 sky130_fd_sc_hs__nand3_1 _07828_ (.A(_02335_),
    .B(\u_dct.n_ptr[2] ),
    .C(\u_dct.n_ptr[1] ),
    .Y(_02343_));
 sky130_fd_sc_hs__nor2_1 _07829_ (.A(_00569_),
    .B(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hs__and2_1 _07830_ (.A(_02343_),
    .B(_00569_),
    .X(_02345_));
 sky130_fd_sc_hs__nor3_1 _07831_ (.A(_02340_),
    .B(_02344_),
    .C(_02345_),
    .Y(_00269_));
 sky130_fd_sc_hs__nor3b_1 _07832_ (.A(_00569_),
    .B(_02341_),
    .C_N(\u_dct.n_ptr[4] ),
    .Y(_02346_));
 sky130_fd_sc_hs__a21oi_1 _07833_ (.A1(_02342_),
    .A2(\u_dct.n_ptr[3] ),
    .B1(\u_dct.n_ptr[4] ),
    .Y(_02347_));
 sky130_fd_sc_hs__nor3_1 _07834_ (.A(_02340_),
    .B(_02346_),
    .C(_02347_),
    .Y(_00270_));
 sky130_fd_sc_hs__and2_1 _07835_ (.A(_02344_),
    .B(\u_dct.n_ptr[4] ),
    .X(_02348_));
 sky130_fd_sc_hs__nor2_1 _07836_ (.A(\u_dct.n_ptr[5] ),
    .B(_02348_),
    .Y(_02349_));
 sky130_fd_sc_hs__and2_1 _07837_ (.A(_02348_),
    .B(\u_dct.n_ptr[5] ),
    .X(_02350_));
 sky130_fd_sc_hs__nor3_1 _07838_ (.A(_02340_),
    .B(_02349_),
    .C(_02350_),
    .Y(_00271_));
 sky130_fd_sc_hs__nor2_1 _07839_ (.A(net3780),
    .B(_02165_),
    .Y(_00272_));
 sky130_fd_sc_hs__nor2_1 _07840_ (.A(_02161_),
    .B(_02156_),
    .Y(_02351_));
 sky130_fd_sc_hs__nor2_1 _07841_ (.A(_02161_),
    .B(_02140_),
    .Y(_02352_));
 sky130_fd_sc_hs__nor2_1 _07842_ (.A(net2991),
    .B(_02352_),
    .Y(_02353_));
 sky130_fd_sc_hs__nor2_1 _07843_ (.A(_02240_),
    .B(_02174_),
    .Y(_02354_));
 sky130_fd_sc_hs__nor2_1 _07844_ (.A(_02161_),
    .B(_02160_),
    .Y(_02355_));
 sky130_fd_sc_hs__nor3_1 _07845_ (.A(_02164_),
    .B(_02354_),
    .C(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hs__nand2_1 _07846_ (.A(_02353_),
    .B(_02356_),
    .Y(_02357_));
 sky130_fd_sc_hs__nor3_1 _07847_ (.A(_02240_),
    .B(\u_fft.power_ptr[0] ),
    .C(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hs__a21oi_1 _07848_ (.A1(\u_fft.power_ptr[0] ),
    .A2(_02357_),
    .B1(_02358_),
    .Y(_02359_));
 sky130_fd_sc_hs__nor2_1 _07849_ (.A(net3780),
    .B(_02359_),
    .Y(_00273_));
 sky130_fd_sc_hs__inv_1 _07850_ (.A(\u_fft.power_ptr[1] ),
    .Y(_02360_));
 sky130_fd_sc_hs__nor2_1 _07851_ (.A(_00202_),
    .B(_02357_),
    .Y(_02361_));
 sky130_fd_sc_hs__o21ai_1 _07852_ (.A1(\u_fft.fft_state[1] ),
    .A2(_02357_),
    .B1(net211),
    .Y(_02362_));
 sky130_fd_sc_hs__a211oi_1 _07853_ (.A1(_02360_),
    .A2(_02357_),
    .B1(_02361_),
    .C1(net2917),
    .Y(_00274_));
 sky130_fd_sc_hs__and3_1 _07854_ (.A(_02353_),
    .B(_00201_),
    .C(_02356_),
    .X(_02363_));
 sky130_fd_sc_hs__nor2_1 _07855_ (.A(\u_fft.power_ptr[2] ),
    .B(_02363_),
    .Y(_02364_));
 sky130_fd_sc_hs__nand2_1 _07856_ (.A(_02363_),
    .B(\u_fft.power_ptr[2] ),
    .Y(_02365_));
 sky130_fd_sc_hs__nor3b_1 _07857_ (.A(net2917),
    .B(_02364_),
    .C_N(_02365_),
    .Y(_00275_));
 sky130_fd_sc_hs__nand3_1 _07858_ (.A(\u_fft.power_ptr[0] ),
    .B(\u_fft.power_ptr[2] ),
    .C(\u_fft.power_ptr[1] ),
    .Y(_02366_));
 sky130_fd_sc_hs__nor2_1 _07859_ (.A(_02366_),
    .B(_02357_),
    .Y(_02367_));
 sky130_fd_sc_hs__xnor2_1 _07860_ (.A(\u_fft.power_ptr[3] ),
    .B(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hs__nor2_1 _07861_ (.A(net2917),
    .B(_02368_),
    .Y(_00276_));
 sky130_fd_sc_hs__clkinv_1 _07862_ (.A(\u_fft.power_ptr[3] ),
    .Y(_02369_));
 sky130_fd_sc_hs__nor2_1 _07863_ (.A(_02369_),
    .B(_02365_),
    .Y(_02370_));
 sky130_fd_sc_hs__nor2_1 _07864_ (.A(\u_fft.power_ptr[4] ),
    .B(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hs__nand2_1 _07865_ (.A(_02370_),
    .B(\u_fft.power_ptr[4] ),
    .Y(_02372_));
 sky130_fd_sc_hs__nor3b_1 _07866_ (.A(net2917),
    .B(_02371_),
    .C_N(_02372_),
    .Y(_00277_));
 sky130_fd_sc_hs__clkinv_1 _07867_ (.A(\u_fft.power_ptr[5] ),
    .Y(_02373_));
 sky130_fd_sc_hs__nand3b_1 _07868_ (.A_N(_02366_),
    .B(\u_fft.power_ptr[3] ),
    .C(\u_fft.power_ptr[4] ),
    .Y(_02374_));
 sky130_fd_sc_hs__nor3_1 _07869_ (.A(_02373_),
    .B(_02374_),
    .C(_02357_),
    .Y(_02375_));
 sky130_fd_sc_hs__nor2_1 _07870_ (.A(_02374_),
    .B(_02357_),
    .Y(_02376_));
 sky130_fd_sc_hs__nor2_1 _07871_ (.A(\u_fft.power_ptr[5] ),
    .B(_02376_),
    .Y(_02377_));
 sky130_fd_sc_hs__nor3_1 _07872_ (.A(net2917),
    .B(_02375_),
    .C(_02377_),
    .Y(_00278_));
 sky130_fd_sc_hs__nor2_1 _07873_ (.A(_02373_),
    .B(_02372_),
    .Y(_02378_));
 sky130_fd_sc_hs__nor2_1 _07874_ (.A(\u_fft.power_ptr[6] ),
    .B(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hs__inv_1 _07875_ (.A(\u_fft.power_ptr[6] ),
    .Y(_02380_));
 sky130_fd_sc_hs__inv_1 _07876_ (.A(_02378_),
    .Y(_02381_));
 sky130_fd_sc_hs__nor2_1 _07877_ (.A(_02380_),
    .B(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hs__nor3_1 _07878_ (.A(net2917),
    .B(_02379_),
    .C(_02382_),
    .Y(_00279_));
 sky130_fd_sc_hs__clkinv_1 _07879_ (.A(\u_fft.power_ptr[7] ),
    .Y(_02383_));
 sky130_fd_sc_hs__nand2_1 _07880_ (.A(_02375_),
    .B(\u_fft.power_ptr[6] ),
    .Y(_02384_));
 sky130_fd_sc_hs__nor2_1 _07881_ (.A(_02383_),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hs__a21oi_1 _07882_ (.A1(_02375_),
    .A2(\u_fft.power_ptr[6] ),
    .B1(\u_fft.power_ptr[7] ),
    .Y(_02386_));
 sky130_fd_sc_hs__nor3_1 _07883_ (.A(net2917),
    .B(_02385_),
    .C(_02386_),
    .Y(_00280_));
 sky130_fd_sc_hs__a21oi_1 _07884_ (.A1(_02382_),
    .A2(\u_fft.power_ptr[7] ),
    .B1(\u_fft.power_ptr[8] ),
    .Y(_02387_));
 sky130_fd_sc_hs__inv_1 _07885_ (.A(\u_fft.power_ptr[8] ),
    .Y(_02388_));
 sky130_fd_sc_hs__nor4_1 _07886_ (.A(_02380_),
    .B(_02383_),
    .C(_02388_),
    .D(_02381_),
    .Y(_02389_));
 sky130_fd_sc_hs__nor3_1 _07887_ (.A(net2917),
    .B(_02387_),
    .C(_02389_),
    .Y(_00281_));
 sky130_fd_sc_hs__a21oi_1 _07888_ (.A1(_02385_),
    .A2(\u_fft.power_ptr[8] ),
    .B1(\u_fft.power_ptr[9] ),
    .Y(_02390_));
 sky130_fd_sc_hs__a31o_1 _07889_ (.A1(_02385_),
    .A2(\u_fft.power_ptr[8] ),
    .A3(\u_fft.power_ptr[9] ),
    .B1(net2917),
    .X(_02391_));
 sky130_fd_sc_hs__nor2_1 _07890_ (.A(_02390_),
    .B(_02391_),
    .Y(_00282_));
 sky130_fd_sc_hs__inv_2 _07891_ (.A(net3338),
    .Y(_02392_));
 sky130_fd_sc_hs__buf_1 place2155 (.A(_05456_),
    .X(net2155));
 sky130_fd_sc_hs__nand2_1 _07893_ (.A(_02392_),
    .B(\u_fft.power_ptr[0] ),
    .Y(_02394_));
 sky130_fd_sc_hs__nand2_1 _07894_ (.A(net3338),
    .B(\u_fft.power_ptr_stage1[0] ),
    .Y(_02395_));
 sky130_fd_sc_hs__a21oi_1 _07895_ (.A1(_02394_),
    .A2(_02395_),
    .B1(net3780),
    .Y(_00283_));
 sky130_fd_sc_hs__o21ai_1 _07896_ (.A1(\u_fft.power_ptr_stage1[1] ),
    .A2(_02392_),
    .B1(net3784),
    .Y(_02396_));
 sky130_fd_sc_hs__a21oi_1 _07897_ (.A1(_02360_),
    .A2(_02392_),
    .B1(_02396_),
    .Y(_00284_));
 sky130_fd_sc_hs__nand2_1 _07898_ (.A(_02392_),
    .B(\u_fft.power_ptr[2] ),
    .Y(_02397_));
 sky130_fd_sc_hs__nand2_1 _07899_ (.A(net3338),
    .B(\u_fft.power_ptr_stage1[2] ),
    .Y(_02398_));
 sky130_fd_sc_hs__a21oi_1 _07900_ (.A1(_02397_),
    .A2(_02398_),
    .B1(_05774_),
    .Y(_00285_));
 sky130_fd_sc_hs__o21ai_1 _07901_ (.A1(\u_fft.power_ptr_stage1[3] ),
    .A2(_02392_),
    .B1(net3784),
    .Y(_02399_));
 sky130_fd_sc_hs__a21oi_1 _07902_ (.A1(_02369_),
    .A2(_02392_),
    .B1(_02399_),
    .Y(_00286_));
 sky130_fd_sc_hs__nand2_1 _07903_ (.A(_02392_),
    .B(\u_fft.power_ptr[4] ),
    .Y(_02400_));
 sky130_fd_sc_hs__nand2_1 _07904_ (.A(net3338),
    .B(\u_fft.power_ptr_stage1[4] ),
    .Y(_02401_));
 sky130_fd_sc_hs__a21oi_1 _07905_ (.A1(_02400_),
    .A2(_02401_),
    .B1(_05774_),
    .Y(_00287_));
 sky130_fd_sc_hs__buf_1 place2173 (.A(_05434_),
    .X(net2173));
 sky130_fd_sc_hs__o21ai_1 _07907_ (.A1(\u_fft.power_ptr_stage1[5] ),
    .A2(_02392_),
    .B1(net3784),
    .Y(_02403_));
 sky130_fd_sc_hs__a21oi_1 _07908_ (.A1(_02373_),
    .A2(_02392_),
    .B1(_02403_),
    .Y(_00288_));
 sky130_fd_sc_hs__o21ai_1 _07909_ (.A1(\u_fft.power_ptr_stage1[6] ),
    .A2(net3300),
    .B1(net211),
    .Y(_02404_));
 sky130_fd_sc_hs__a21oi_1 _07910_ (.A1(_02380_),
    .A2(net3300),
    .B1(_02404_),
    .Y(_00289_));
 sky130_fd_sc_hs__o21ai_1 _07911_ (.A1(\u_fft.power_ptr_stage1[7] ),
    .A2(net3300),
    .B1(net211),
    .Y(_02405_));
 sky130_fd_sc_hs__a21oi_1 _07912_ (.A1(_02383_),
    .A2(net3300),
    .B1(_02405_),
    .Y(_00290_));
 sky130_fd_sc_hs__o21ai_1 _07913_ (.A1(\u_fft.power_ptr_stage1[8] ),
    .A2(net3300),
    .B1(net211),
    .Y(_02406_));
 sky130_fd_sc_hs__a21oi_1 _07914_ (.A1(_02388_),
    .A2(net3300),
    .B1(_02406_),
    .Y(_00291_));
 sky130_fd_sc_hs__nand2_1 _07915_ (.A(net3300),
    .B(\u_fft.power_ptr[9] ),
    .Y(_02407_));
 sky130_fd_sc_hs__nand2_1 _07916_ (.A(net3338),
    .B(\u_fft.power_ptr_stage1[9] ),
    .Y(_02408_));
 sky130_fd_sc_hs__a21oi_1 _07917_ (.A1(_02407_),
    .A2(_02408_),
    .B1(net3781),
    .Y(_00292_));
 sky130_fd_sc_hs__buf_2 place2154 (.A(_03489_),
    .X(net2154));
 sky130_fd_sc_hs__nand2_1 _07919_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage1[0] ),
    .Y(_02410_));
 sky130_fd_sc_hs__nand2_1 _07920_ (.A(net3338),
    .B(\u_fft.power_ptr_stage2[0] ),
    .Y(_02411_));
 sky130_fd_sc_hs__a21oi_1 _07921_ (.A1(_02410_),
    .A2(_02411_),
    .B1(net3780),
    .Y(_00293_));
 sky130_fd_sc_hs__nand2_1 _07922_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage1[1] ),
    .Y(_02412_));
 sky130_fd_sc_hs__nand2_1 _07923_ (.A(net3338),
    .B(\u_fft.power_ptr_stage2[1] ),
    .Y(_02413_));
 sky130_fd_sc_hs__a21oi_1 _07924_ (.A1(_02412_),
    .A2(_02413_),
    .B1(net3780),
    .Y(_00294_));
 sky130_fd_sc_hs__nand2_1 _07925_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage1[2] ),
    .Y(_02414_));
 sky130_fd_sc_hs__nand2_1 _07926_ (.A(net3338),
    .B(\u_fft.power_ptr_stage2[2] ),
    .Y(_02415_));
 sky130_fd_sc_hs__a21oi_1 _07927_ (.A1(_02414_),
    .A2(_02415_),
    .B1(_05774_),
    .Y(_00295_));
 sky130_fd_sc_hs__nand2_1 _07928_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage1[3] ),
    .Y(_02416_));
 sky130_fd_sc_hs__nand2_1 _07929_ (.A(net3338),
    .B(\u_fft.power_ptr_stage2[3] ),
    .Y(_02417_));
 sky130_fd_sc_hs__a21oi_1 _07930_ (.A1(_02416_),
    .A2(_02417_),
    .B1(_05774_),
    .Y(_00296_));
 sky130_fd_sc_hs__nand2_1 _07931_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage1[4] ),
    .Y(_02418_));
 sky130_fd_sc_hs__nand2_1 _07932_ (.A(net3338),
    .B(\u_fft.power_ptr_stage2[4] ),
    .Y(_02419_));
 sky130_fd_sc_hs__buf_1 place2152 (.A(_04561_),
    .X(net2152));
 sky130_fd_sc_hs__a21oi_1 _07934_ (.A1(_02418_),
    .A2(_02419_),
    .B1(_05774_),
    .Y(_00297_));
 sky130_fd_sc_hs__nand2_1 _07935_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage1[5] ),
    .Y(_02421_));
 sky130_fd_sc_hs__buf_1 place2151 (.A(_05461_),
    .X(net2151));
 sky130_fd_sc_hs__nand2_1 _07937_ (.A(net3338),
    .B(\u_fft.power_ptr_stage2[5] ),
    .Y(_02423_));
 sky130_fd_sc_hs__a21oi_1 _07938_ (.A1(_02421_),
    .A2(_02423_),
    .B1(_05774_),
    .Y(_00298_));
 sky130_fd_sc_hs__nand2_1 _07939_ (.A(net3300),
    .B(\u_fft.power_ptr_stage1[6] ),
    .Y(_02424_));
 sky130_fd_sc_hs__nand2_1 _07940_ (.A(net3338),
    .B(\u_fft.power_ptr_stage2[6] ),
    .Y(_02425_));
 sky130_fd_sc_hs__a21oi_1 _07941_ (.A1(_02424_),
    .A2(_02425_),
    .B1(net3781),
    .Y(_00299_));
 sky130_fd_sc_hs__nand2_1 _07942_ (.A(net3300),
    .B(\u_fft.power_ptr_stage1[7] ),
    .Y(_02426_));
 sky130_fd_sc_hs__nand2_1 _07943_ (.A(net3338),
    .B(\u_fft.power_ptr_stage2[7] ),
    .Y(_02427_));
 sky130_fd_sc_hs__a21oi_1 _07944_ (.A1(_02426_),
    .A2(_02427_),
    .B1(_05774_),
    .Y(_00300_));
 sky130_fd_sc_hs__nand2_1 _07945_ (.A(net3300),
    .B(\u_fft.power_ptr_stage1[8] ),
    .Y(_02428_));
 sky130_fd_sc_hs__nand2_1 _07946_ (.A(net3338),
    .B(\u_fft.power_ptr_stage2[8] ),
    .Y(_02429_));
 sky130_fd_sc_hs__a21oi_1 _07947_ (.A1(_02428_),
    .A2(_02429_),
    .B1(net3781),
    .Y(_00301_));
 sky130_fd_sc_hs__nand2_1 _07948_ (.A(net3300),
    .B(\u_fft.power_ptr_stage1[9] ),
    .Y(_02430_));
 sky130_fd_sc_hs__nand2_1 _07949_ (.A(net3338),
    .B(\u_fft.power_ptr_stage2[9] ),
    .Y(_02431_));
 sky130_fd_sc_hs__a21oi_1 _07950_ (.A1(_02430_),
    .A2(_02431_),
    .B1(net3781),
    .Y(_00302_));
 sky130_fd_sc_hs__buf_1 place2149 (.A(_05476_),
    .X(net2149));
 sky130_fd_sc_hs__nand2_1 _07952_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage2[0] ),
    .Y(_02433_));
 sky130_fd_sc_hs__nand2_1 _07953_ (.A(net3338),
    .B(\u_fft.power_ptr_stage3[0] ),
    .Y(_02434_));
 sky130_fd_sc_hs__a21oi_1 _07954_ (.A1(_02433_),
    .A2(_02434_),
    .B1(net3780),
    .Y(_00303_));
 sky130_fd_sc_hs__nand2_1 _07955_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage2[1] ),
    .Y(_02435_));
 sky130_fd_sc_hs__nand2_1 _07956_ (.A(net3338),
    .B(\u_fft.power_ptr_stage3[1] ),
    .Y(_02436_));
 sky130_fd_sc_hs__a21oi_1 _07957_ (.A1(_02435_),
    .A2(_02436_),
    .B1(net3780),
    .Y(_00304_));
 sky130_fd_sc_hs__nand2_1 _07958_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage2[2] ),
    .Y(_02437_));
 sky130_fd_sc_hs__nand2_1 _07959_ (.A(net3338),
    .B(\u_fft.power_ptr_stage3[2] ),
    .Y(_02438_));
 sky130_fd_sc_hs__a21oi_1 _07960_ (.A1(_02437_),
    .A2(_02438_),
    .B1(_05774_),
    .Y(_00305_));
 sky130_fd_sc_hs__nand2_1 _07961_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage2[3] ),
    .Y(_02439_));
 sky130_fd_sc_hs__nand2_1 _07962_ (.A(net3338),
    .B(\u_fft.power_ptr_stage3[3] ),
    .Y(_02440_));
 sky130_fd_sc_hs__a21oi_1 _07963_ (.A1(_02439_),
    .A2(_02440_),
    .B1(_05774_),
    .Y(_00306_));
 sky130_fd_sc_hs__nand2_1 _07964_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage2[4] ),
    .Y(_02441_));
 sky130_fd_sc_hs__nand2_1 _07965_ (.A(net3338),
    .B(\u_fft.power_ptr_stage3[4] ),
    .Y(_02442_));
 sky130_fd_sc_hs__buf_1 place2148 (.A(_05484_),
    .X(net2148));
 sky130_fd_sc_hs__a21oi_1 _07967_ (.A1(_02441_),
    .A2(_02442_),
    .B1(_05774_),
    .Y(_00307_));
 sky130_fd_sc_hs__nand2_1 _07968_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage2[5] ),
    .Y(_02444_));
 sky130_fd_sc_hs__buf_1 place2147 (.A(_01718_),
    .X(net2147));
 sky130_fd_sc_hs__nand2_1 _07970_ (.A(net3338),
    .B(\u_fft.power_ptr_stage3[5] ),
    .Y(_02446_));
 sky130_fd_sc_hs__a21oi_1 _07971_ (.A1(_02444_),
    .A2(_02446_),
    .B1(_05774_),
    .Y(_00308_));
 sky130_fd_sc_hs__nand2_1 _07972_ (.A(net3300),
    .B(\u_fft.power_ptr_stage2[6] ),
    .Y(_02447_));
 sky130_fd_sc_hs__nand2_1 _07973_ (.A(net3338),
    .B(\u_fft.power_ptr_stage3[6] ),
    .Y(_02448_));
 sky130_fd_sc_hs__a21oi_1 _07974_ (.A1(_02447_),
    .A2(_02448_),
    .B1(net3781),
    .Y(_00309_));
 sky130_fd_sc_hs__nand2_1 _07975_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage2[7] ),
    .Y(_02449_));
 sky130_fd_sc_hs__nand2_1 _07976_ (.A(net3338),
    .B(\u_fft.power_ptr_stage3[7] ),
    .Y(_02450_));
 sky130_fd_sc_hs__a21oi_1 _07977_ (.A1(_02449_),
    .A2(_02450_),
    .B1(_05774_),
    .Y(_00310_));
 sky130_fd_sc_hs__nand2_1 _07978_ (.A(net3300),
    .B(\u_fft.power_ptr_stage2[8] ),
    .Y(_02451_));
 sky130_fd_sc_hs__nand2_1 _07979_ (.A(net3338),
    .B(\u_fft.power_ptr_stage3[8] ),
    .Y(_02452_));
 sky130_fd_sc_hs__a21oi_1 _07980_ (.A1(_02451_),
    .A2(_02452_),
    .B1(net3781),
    .Y(_00311_));
 sky130_fd_sc_hs__nand2_1 _07981_ (.A(net3300),
    .B(\u_fft.power_ptr_stage2[9] ),
    .Y(_02453_));
 sky130_fd_sc_hs__nand2_1 _07982_ (.A(net3338),
    .B(\u_fft.power_ptr_stage3[9] ),
    .Y(_02454_));
 sky130_fd_sc_hs__a21oi_1 _07983_ (.A1(_02453_),
    .A2(_02454_),
    .B1(net3781),
    .Y(_00312_));
 sky130_fd_sc_hs__buf_1 place2146 (.A(_03483_),
    .X(net2146));
 sky130_fd_sc_hs__nand2_1 _07985_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage3[0] ),
    .Y(_02456_));
 sky130_fd_sc_hs__nand2_1 _07986_ (.A(net3338),
    .B(\fft_ptr[0] ),
    .Y(_02457_));
 sky130_fd_sc_hs__a21oi_1 _07987_ (.A1(_02456_),
    .A2(_02457_),
    .B1(_05774_),
    .Y(_00313_));
 sky130_fd_sc_hs__nand2_1 _07988_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage3[1] ),
    .Y(_02458_));
 sky130_fd_sc_hs__nand2_1 _07989_ (.A(net3338),
    .B(\fft_ptr[1] ),
    .Y(_02459_));
 sky130_fd_sc_hs__a21oi_1 _07990_ (.A1(_02458_),
    .A2(_02459_),
    .B1(_05774_),
    .Y(_00314_));
 sky130_fd_sc_hs__nand2_1 _07991_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage3[2] ),
    .Y(_02460_));
 sky130_fd_sc_hs__nand2_1 _07992_ (.A(net3338),
    .B(\fft_ptr[2] ),
    .Y(_02461_));
 sky130_fd_sc_hs__a21oi_1 _07993_ (.A1(_02460_),
    .A2(_02461_),
    .B1(_05774_),
    .Y(_00315_));
 sky130_fd_sc_hs__nand2_1 _07994_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage3[3] ),
    .Y(_02462_));
 sky130_fd_sc_hs__nand2_1 _07995_ (.A(net3338),
    .B(\fft_ptr[3] ),
    .Y(_02463_));
 sky130_fd_sc_hs__a21oi_1 _07996_ (.A1(_02462_),
    .A2(_02463_),
    .B1(_05774_),
    .Y(_00316_));
 sky130_fd_sc_hs__nand2_1 _07997_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage3[4] ),
    .Y(_02464_));
 sky130_fd_sc_hs__nand2_1 _07998_ (.A(net3338),
    .B(\fft_ptr[4] ),
    .Y(_02465_));
 sky130_fd_sc_hs__buf_1 place2145 (.A(_04558_),
    .X(net2145));
 sky130_fd_sc_hs__a21oi_1 _08000_ (.A1(_02464_),
    .A2(_02465_),
    .B1(_05774_),
    .Y(_00317_));
 sky130_fd_sc_hs__nand2_1 _08001_ (.A(_02392_),
    .B(\u_fft.power_ptr_stage3[5] ),
    .Y(_02467_));
 sky130_fd_sc_hs__nand2_1 _08002_ (.A(net3338),
    .B(\fft_ptr[5] ),
    .Y(_02468_));
 sky130_fd_sc_hs__a21oi_1 _08003_ (.A1(_02467_),
    .A2(_02468_),
    .B1(_05774_),
    .Y(_00318_));
 sky130_fd_sc_hs__nand2_1 _08004_ (.A(net3300),
    .B(\u_fft.power_ptr_stage3[6] ),
    .Y(_02469_));
 sky130_fd_sc_hs__nand2_1 _08005_ (.A(net3338),
    .B(\fft_ptr[6] ),
    .Y(_02470_));
 sky130_fd_sc_hs__a21oi_1 _08006_ (.A1(_02469_),
    .A2(_02470_),
    .B1(net3781),
    .Y(_00319_));
 sky130_fd_sc_hs__nand2_1 _08007_ (.A(net3300),
    .B(\u_fft.power_ptr_stage3[7] ),
    .Y(_02471_));
 sky130_fd_sc_hs__nand2_1 _08008_ (.A(net3338),
    .B(\fft_ptr[7] ),
    .Y(_02472_));
 sky130_fd_sc_hs__a21oi_1 _08009_ (.A1(_02471_),
    .A2(_02472_),
    .B1(net3781),
    .Y(_00320_));
 sky130_fd_sc_hs__nand2_1 _08010_ (.A(net3300),
    .B(\u_fft.power_ptr_stage3[8] ),
    .Y(_02473_));
 sky130_fd_sc_hs__nand2_1 _08011_ (.A(net3338),
    .B(\fft_ptr[8] ),
    .Y(_02474_));
 sky130_fd_sc_hs__a21oi_1 _08012_ (.A1(_02473_),
    .A2(_02474_),
    .B1(net3781),
    .Y(_00321_));
 sky130_fd_sc_hs__nand2_1 _08013_ (.A(net3300),
    .B(\u_fft.power_ptr_stage3[9] ),
    .Y(_02475_));
 sky130_fd_sc_hs__nand2_1 _08014_ (.A(net3338),
    .B(\u_fft.power_ptr_stage4[9] ),
    .Y(_02476_));
 sky130_fd_sc_hs__a21oi_1 _08015_ (.A1(_02475_),
    .A2(_02476_),
    .B1(net3781),
    .Y(_00322_));
 sky130_fd_sc_hs__a21oi_1 _08016_ (.A1(_02161_),
    .A2(_02163_),
    .B1(_02164_),
    .Y(_02477_));
 sky130_fd_sc_hs__inv_2 _08017_ (.A(_02477_),
    .Y(_02478_));
 sky130_fd_sc_hs__nor2_1 _08018_ (.A(_02478_),
    .B(_02352_),
    .Y(_02479_));
 sky130_fd_sc_hs__nor2_1 _08019_ (.A(_02167_),
    .B(_02351_),
    .Y(_02480_));
 sky130_fd_sc_hs__nand2_1 _08020_ (.A(_02479_),
    .B(_02480_),
    .Y(_02481_));
 sky130_fd_sc_hs__buf_1 place2144 (.A(_04563_),
    .X(net2144));
 sky130_fd_sc_hs__inv_2 _08022_ (.A(net2941),
    .Y(_02483_));
 sky130_fd_sc_hs__buf_2 place2143 (.A(_05475_),
    .X(net2143));
 sky130_fd_sc_hs__nor2_1 _08024_ (.A(\u_fft.sched[20] ),
    .B(_02483_),
    .Y(_02485_));
 sky130_fd_sc_hs__inv_1 _08025_ (.A(_00171_),
    .Y(_02486_));
 sky130_fd_sc_hs__nor2_1 _08026_ (.A(\u_fft.sched[42] ),
    .B(_02486_),
    .Y(_02487_));
 sky130_fd_sc_hs__nor2_1 _08027_ (.A(_02161_),
    .B(_02481_),
    .Y(_02488_));
 sky130_fd_sc_hs__inv_2 _08028_ (.A(_02488_),
    .Y(_02489_));
 sky130_fd_sc_hs__a21oi_1 _08029_ (.A1(_02159_),
    .A2(_02487_),
    .B1(_02489_),
    .Y(_02490_));
 sky130_fd_sc_hs__o21ai_1 _08030_ (.A1(_02485_),
    .A2(_02490_),
    .B1(net211),
    .Y(_00323_));
 sky130_fd_sc_hs__buf_1 place2142 (.A(_05487_),
    .X(net2142));
 sky130_fd_sc_hs__nand2_1 _08032_ (.A(_02159_),
    .B(\u_fft.fft_state[2] ),
    .Y(_02492_));
 sky130_fd_sc_hs__inv_1 _08033_ (.A(_02492_),
    .Y(_02493_));
 sky130_fd_sc_hs__a31oi_1 _08034_ (.A1(_00176_),
    .A2(_00174_),
    .A3(_02493_),
    .B1(_02481_),
    .Y(_02494_));
 sky130_fd_sc_hs__a211oi_1 _08035_ (.A1(_02481_),
    .A2(_00054_),
    .B1(net3780),
    .C1(_02494_),
    .Y(_00324_));
 sky130_fd_sc_hs__nor2_1 _08036_ (.A(\u_fft.sched[22] ),
    .B(_02483_),
    .Y(_02495_));
 sky130_fd_sc_hs__buf_1 place2141 (.A(_01716_),
    .X(net2141));
 sky130_fd_sc_hs__a31oi_1 _08038_ (.A1(_00176_),
    .A2(_00173_),
    .A3(_02493_),
    .B1(_02481_),
    .Y(_02497_));
 sky130_fd_sc_hs__nor3_1 _08039_ (.A(net3780),
    .B(_02495_),
    .C(_02497_),
    .Y(_00325_));
 sky130_fd_sc_hs__a21oi_1 _08040_ (.A1(_00177_),
    .A2(_02493_),
    .B1(_02481_),
    .Y(_02498_));
 sky130_fd_sc_hs__a211oi_1 _08041_ (.A1(_05781_),
    .A2(_02481_),
    .B1(net3780),
    .C1(_02498_),
    .Y(_00326_));
 sky130_fd_sc_hs__nor2_1 _08042_ (.A(_00176_),
    .B(_02492_),
    .Y(_02499_));
 sky130_fd_sc_hs__a21oi_1 _08043_ (.A1(_00171_),
    .A2(_02499_),
    .B1(_02481_),
    .Y(_02500_));
 sky130_fd_sc_hs__a211oi_1 _08044_ (.A1(_05780_),
    .A2(_02481_),
    .B1(net3780),
    .C1(_02500_),
    .Y(_00327_));
 sky130_fd_sc_hs__a21oi_1 _08045_ (.A1(_00174_),
    .A2(_02499_),
    .B1(_02481_),
    .Y(_02501_));
 sky130_fd_sc_hs__nor2_1 _08046_ (.A(\u_fft.sched[25] ),
    .B(_02483_),
    .Y(_02502_));
 sky130_fd_sc_hs__nor3_1 _08047_ (.A(net3780),
    .B(_02501_),
    .C(_02502_),
    .Y(_00328_));
 sky130_fd_sc_hs__a21oi_1 _08048_ (.A1(_00173_),
    .A2(_02499_),
    .B1(_02481_),
    .Y(_02503_));
 sky130_fd_sc_hs__nor2_1 _08049_ (.A(\u_fft.sched[26] ),
    .B(_02483_),
    .Y(_02504_));
 sky130_fd_sc_hs__nor3_1 _08050_ (.A(net3780),
    .B(_02503_),
    .C(_02504_),
    .Y(_00329_));
 sky130_fd_sc_hs__a21oi_1 _08051_ (.A1(_00179_),
    .A2(_02493_),
    .B1(_02481_),
    .Y(_02505_));
 sky130_fd_sc_hs__nor2_1 _08052_ (.A(\u_fft.sched[1] ),
    .B(_02483_),
    .Y(_02506_));
 sky130_fd_sc_hs__nor3_1 _08053_ (.A(net3780),
    .B(_02505_),
    .C(_02506_),
    .Y(_00330_));
 sky130_fd_sc_hs__inv_1 _08054_ (.A(\u_fft.sched[43] ),
    .Y(_02507_));
 sky130_fd_sc_hs__nor3_1 _08055_ (.A(\u_fft.sched[44] ),
    .B(_02161_),
    .C(_02507_),
    .Y(_02508_));
 sky130_fd_sc_hs__a21oi_1 _08056_ (.A1(_02487_),
    .A2(_02508_),
    .B1(_02481_),
    .Y(_02509_));
 sky130_fd_sc_hs__nor2_1 _08057_ (.A(\u_fft.sched[0] ),
    .B(_02483_),
    .Y(_02510_));
 sky130_fd_sc_hs__nor3_1 _08058_ (.A(net3780),
    .B(_02509_),
    .C(_02510_),
    .Y(_00331_));
 sky130_fd_sc_hs__nor2_1 _08059_ (.A(\u_fft.sched[29] ),
    .B(_02483_),
    .Y(_02511_));
 sky130_fd_sc_hs__a31oi_1 _08060_ (.A1(_00176_),
    .A2(_00174_),
    .A3(_02508_),
    .B1(_02481_),
    .Y(_02512_));
 sky130_fd_sc_hs__nor3_1 _08061_ (.A(net3780),
    .B(_02511_),
    .C(_02512_),
    .Y(_00332_));
 sky130_fd_sc_hs__buf_4 place2140 (.A(_03473_),
    .X(net2140));
 sky130_fd_sc_hs__inv_1 _08063_ (.A(_00178_),
    .Y(_02514_));
 sky130_fd_sc_hs__nand3_1 _08064_ (.A(\u_fft.sched[43] ),
    .B(\u_fft.sched[42] ),
    .C(_00175_),
    .Y(_02515_));
 sky130_fd_sc_hs__xnor2_1 _08065_ (.A(_02158_),
    .B(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hs__inv_1 _08066_ (.A(_02516_),
    .Y(_02517_));
 sky130_fd_sc_hs__nor2_1 _08067_ (.A(_00176_),
    .B(_00170_),
    .Y(_02518_));
 sky130_fd_sc_hs__a31oi_1 _08068_ (.A1(_02518_),
    .A2(\u_fft.sched[44] ),
    .A3(\u_fft.sched[43] ),
    .B1(_00169_),
    .Y(_02519_));
 sky130_fd_sc_hs__inv_2 _08069_ (.A(_02519_),
    .Y(_02520_));
 sky130_fd_sc_hs__nor4_1 _08070_ (.A(_02514_),
    .B(_00172_),
    .C(_02517_),
    .D(_02520_),
    .Y(_02521_));
 sky130_fd_sc_hs__nand2_1 _08071_ (.A(_02518_),
    .B(\u_fft.sched[40] ),
    .Y(_02522_));
 sky130_fd_sc_hs__xnor2_1 _08072_ (.A(_02507_),
    .B(_02522_),
    .Y(_02523_));
 sky130_fd_sc_hs__a31oi_1 _08073_ (.A1(\u_fft.fft_state[2] ),
    .A2(_02521_),
    .A3(_02523_),
    .B1(net2941),
    .Y(_02524_));
 sky130_fd_sc_hs__a211oi_1 _08074_ (.A1(net2941),
    .A2(_00082_),
    .B1(net3780),
    .C1(_02524_),
    .Y(_00333_));
 sky130_fd_sc_hs__nor2_1 _08075_ (.A(\u_fft.sched[31] ),
    .B(_02483_),
    .Y(_02525_));
 sky130_fd_sc_hs__nor3_1 _08076_ (.A(_02514_),
    .B(_02486_),
    .C(_02517_),
    .Y(_02526_));
 sky130_fd_sc_hs__a21oi_1 _08077_ (.A1(_02523_),
    .A2(_02526_),
    .B1(_02489_),
    .Y(_02527_));
 sky130_fd_sc_hs__o21ai_1 _08078_ (.A1(_02525_),
    .A2(_02527_),
    .B1(net211),
    .Y(_00334_));
 sky130_fd_sc_hs__nor2_1 _08079_ (.A(_02161_),
    .B(_02514_),
    .Y(_02528_));
 sky130_fd_sc_hs__nand2_1 _08080_ (.A(_02523_),
    .B(_02516_),
    .Y(_02529_));
 sky130_fd_sc_hs__nor3b_1 _08081_ (.A(_02529_),
    .B(_02520_),
    .C_N(_00172_),
    .Y(_02530_));
 sky130_fd_sc_hs__a21oi_1 _08082_ (.A1(_02528_),
    .A2(_02530_),
    .B1(net2941),
    .Y(_02531_));
 sky130_fd_sc_hs__nor2_1 _08083_ (.A(\u_fft.sched[32] ),
    .B(_02483_),
    .Y(_02532_));
 sky130_fd_sc_hs__nor3_1 _08084_ (.A(net3780),
    .B(_02531_),
    .C(_02532_),
    .Y(_00335_));
 sky130_fd_sc_hs__nand2_1 _08085_ (.A(_02528_),
    .B(_00173_),
    .Y(_02533_));
 sky130_fd_sc_hs__nor3_1 _08086_ (.A(_02529_),
    .B(_02533_),
    .C(net2941),
    .Y(_02534_));
 sky130_fd_sc_hs__a21oi_1 _08087_ (.A1(\u_fft.sched[33] ),
    .A2(net2941),
    .B1(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hs__nor2_1 _08088_ (.A(net3780),
    .B(_02535_),
    .Y(_00336_));
 sky130_fd_sc_hs__nor2_1 _08089_ (.A(_00172_),
    .B(_02520_),
    .Y(_02536_));
 sky130_fd_sc_hs__nand2_1 _08090_ (.A(_02523_),
    .B(\u_fft.fft_state[2] ),
    .Y(_02537_));
 sky130_fd_sc_hs__nor3_1 _08091_ (.A(_00178_),
    .B(_02517_),
    .C(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hs__a21oi_1 _08092_ (.A1(_02536_),
    .A2(_02538_),
    .B1(net2941),
    .Y(_02539_));
 sky130_fd_sc_hs__nor2_1 _08093_ (.A(\u_fft.sched[34] ),
    .B(_02483_),
    .Y(_02540_));
 sky130_fd_sc_hs__nor3_1 _08094_ (.A(net3780),
    .B(_02539_),
    .C(_02540_),
    .Y(_00337_));
 sky130_fd_sc_hs__a21oi_1 _08095_ (.A1(_00171_),
    .A2(_02538_),
    .B1(net2941),
    .Y(_02541_));
 sky130_fd_sc_hs__nor2_1 _08096_ (.A(\u_fft.sched[35] ),
    .B(_02483_),
    .Y(_02542_));
 sky130_fd_sc_hs__nor3_1 _08097_ (.A(net3780),
    .B(_02541_),
    .C(_02542_),
    .Y(_00338_));
 sky130_fd_sc_hs__nor2_1 _08098_ (.A(_00178_),
    .B(_02489_),
    .Y(_02543_));
 sky130_fd_sc_hs__nand2_1 _08099_ (.A(_02543_),
    .B(_02530_),
    .Y(_02544_));
 sky130_fd_sc_hs__nand2_1 _08100_ (.A(net2941),
    .B(\u_fft.sched[36] ),
    .Y(_02545_));
 sky130_fd_sc_hs__a21oi_1 _08101_ (.A1(_02544_),
    .A2(_02545_),
    .B1(net3780),
    .Y(_00339_));
 sky130_fd_sc_hs__a21oi_1 _08102_ (.A1(_00173_),
    .A2(_02538_),
    .B1(net2941),
    .Y(_02546_));
 sky130_fd_sc_hs__a211oi_1 _08103_ (.A1(_05795_),
    .A2(net2941),
    .B1(net3780),
    .C1(_02546_),
    .Y(_00340_));
 sky130_fd_sc_hs__nor2_1 _08104_ (.A(_02523_),
    .B(_02489_),
    .Y(_02547_));
 sky130_fd_sc_hs__nand2_1 _08105_ (.A(_02547_),
    .B(_02521_),
    .Y(_02548_));
 sky130_fd_sc_hs__nand2_1 _08106_ (.A(net2941),
    .B(\u_fft.sched[38] ),
    .Y(_02549_));
 sky130_fd_sc_hs__a21oi_1 _08107_ (.A1(_02548_),
    .A2(_02549_),
    .B1(net3780),
    .Y(_00341_));
 sky130_fd_sc_hs__nand2_1 _08108_ (.A(_02547_),
    .B(_02526_),
    .Y(_02550_));
 sky130_fd_sc_hs__nand2_1 _08109_ (.A(net2941),
    .B(\u_fft.sched[39] ),
    .Y(_02551_));
 sky130_fd_sc_hs__a21oi_1 _08110_ (.A1(_02550_),
    .A2(_02551_),
    .B1(net3780),
    .Y(_00342_));
 sky130_fd_sc_hs__buf_1 place2137 (.A(_03495_),
    .X(net2137));
 sky130_fd_sc_hs__a21oi_1 _08112_ (.A1(_02483_),
    .A2(_00169_),
    .B1(net3780),
    .Y(_02553_));
 sky130_fd_sc_hs__o21ai_1 _08113_ (.A1(_00169_),
    .A2(_02488_),
    .B1(_02553_),
    .Y(_00343_));
 sky130_fd_sc_hs__nand2_1 _08114_ (.A(_02488_),
    .B(_00172_),
    .Y(_02554_));
 sky130_fd_sc_hs__nand2_1 _08115_ (.A(net2941),
    .B(\u_fft.sched[41] ),
    .Y(_02555_));
 sky130_fd_sc_hs__a21oi_1 _08116_ (.A1(_02554_),
    .A2(_02555_),
    .B1(net3780),
    .Y(_00344_));
 sky130_fd_sc_hs__a21oi_1 _08117_ (.A1(\u_fft.sched[42] ),
    .A2(net2941),
    .B1(_02543_),
    .Y(_02556_));
 sky130_fd_sc_hs__nor2_1 _08118_ (.A(net3780),
    .B(_02556_),
    .Y(_00345_));
 sky130_fd_sc_hs__a21oi_1 _08119_ (.A1(\u_fft.sched[43] ),
    .A2(net2941),
    .B1(_02547_),
    .Y(_02557_));
 sky130_fd_sc_hs__nor2_1 _08120_ (.A(net3780),
    .B(_02557_),
    .Y(_00346_));
 sky130_fd_sc_hs__nor3_1 _08121_ (.A(net3780),
    .B(_02158_),
    .C(_02483_),
    .Y(_00347_));
 sky130_fd_sc_hs__xnor2_1 _08122_ (.A(\u_fft.sched[45] ),
    .B(_02477_),
    .Y(_02558_));
 sky130_fd_sc_hs__inv_2 _08123_ (.A(net2960),
    .Y(_02559_));
 sky130_fd_sc_hs__nand2_1 _08124_ (.A(_02559_),
    .B(net211),
    .Y(_02560_));
 sky130_fd_sc_hs__nor2_1 _08125_ (.A(_02558_),
    .B(_02560_),
    .Y(_00348_));
 sky130_fd_sc_hs__nand3_1 _08126_ (.A(_02352_),
    .B(_00181_),
    .C(_02477_),
    .Y(_02561_));
 sky130_fd_sc_hs__nand2_1 _08127_ (.A(_02478_),
    .B(\u_fft.sched[46] ),
    .Y(_02562_));
 sky130_fd_sc_hs__buf_1 place2134 (.A(_04579_),
    .X(net2134));
 sky130_fd_sc_hs__a21oi_1 _08129_ (.A1(_02561_),
    .A2(_02562_),
    .B1(net3780),
    .Y(_00349_));
 sky130_fd_sc_hs__inv_1 _08130_ (.A(\u_fft.sched[47] ),
    .Y(_02564_));
 sky130_fd_sc_hs__nand2_1 _08131_ (.A(_02477_),
    .B(_00180_),
    .Y(_02565_));
 sky130_fd_sc_hs__xnor2_1 _08132_ (.A(_02564_),
    .B(_02565_),
    .Y(_02566_));
 sky130_fd_sc_hs__nor2_1 _08133_ (.A(_02566_),
    .B(_02560_),
    .Y(_00350_));
 sky130_fd_sc_hs__and2_1 _08134_ (.A(\u_fft.sched[47] ),
    .B(\u_fft.sched[46] ),
    .X(_02567_));
 sky130_fd_sc_hs__and2_1 _08135_ (.A(_02567_),
    .B(\u_fft.sched[45] ),
    .X(_02568_));
 sky130_fd_sc_hs__nand2_1 _08136_ (.A(_02477_),
    .B(_02568_),
    .Y(_02569_));
 sky130_fd_sc_hs__xor2_1 _08137_ (.A(\u_fft.sched[48] ),
    .B(_02569_),
    .X(_02570_));
 sky130_fd_sc_hs__nor2_1 _08138_ (.A(_02570_),
    .B(_02560_),
    .Y(_00351_));
 sky130_fd_sc_hs__nand3_1 _08139_ (.A(\u_fft.sched[47] ),
    .B(_00180_),
    .C(\u_fft.sched[48] ),
    .Y(_02571_));
 sky130_fd_sc_hs__nor2_1 _08140_ (.A(_02571_),
    .B(_02478_),
    .Y(_02572_));
 sky130_fd_sc_hs__xnor2_1 _08141_ (.A(\u_fft.sched[49] ),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hs__nor2_1 _08142_ (.A(_02573_),
    .B(_02560_),
    .Y(_00352_));
 sky130_fd_sc_hs__nand3_1 _08143_ (.A(_02568_),
    .B(\u_fft.sched[49] ),
    .C(\u_fft.sched[48] ),
    .Y(_02574_));
 sky130_fd_sc_hs__nor2_1 _08144_ (.A(_02574_),
    .B(_02478_),
    .Y(_02575_));
 sky130_fd_sc_hs__nor2_1 _08145_ (.A(\u_fft.sched[50] ),
    .B(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hs__nand2_1 _08146_ (.A(_02575_),
    .B(\u_fft.sched[50] ),
    .Y(_02577_));
 sky130_fd_sc_hs__nor3b_1 _08147_ (.A(_02576_),
    .B(_02560_),
    .C_N(_02577_),
    .Y(_00353_));
 sky130_fd_sc_hs__inv_2 _08148_ (.A(\u_fft.sched[51] ),
    .Y(_02578_));
 sky130_fd_sc_hs__nand3_1 _08149_ (.A(_02572_),
    .B(\u_fft.sched[50] ),
    .C(\u_fft.sched[49] ),
    .Y(_02579_));
 sky130_fd_sc_hs__nor2_1 _08150_ (.A(_02578_),
    .B(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hs__and2_1 _08151_ (.A(_02579_),
    .B(_02578_),
    .X(_02581_));
 sky130_fd_sc_hs__nor3_1 _08152_ (.A(_02580_),
    .B(_02581_),
    .C(_02560_),
    .Y(_00354_));
 sky130_fd_sc_hs__nor2_1 _08153_ (.A(_02578_),
    .B(_02577_),
    .Y(_02582_));
 sky130_fd_sc_hs__nor2_1 _08154_ (.A(\u_fft.sched[52] ),
    .B(_02582_),
    .Y(_02583_));
 sky130_fd_sc_hs__nand2_1 _08155_ (.A(_02582_),
    .B(\u_fft.sched[52] ),
    .Y(_02584_));
 sky130_fd_sc_hs__nor3b_1 _08156_ (.A(_02583_),
    .B(_02560_),
    .C_N(_02584_),
    .Y(_00355_));
 sky130_fd_sc_hs__inv_2 _08157_ (.A(\u_fft.sched[53] ),
    .Y(_02585_));
 sky130_fd_sc_hs__nand2_1 _08158_ (.A(_02580_),
    .B(\u_fft.sched[52] ),
    .Y(_02586_));
 sky130_fd_sc_hs__xnor2_1 _08159_ (.A(_02585_),
    .B(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hs__nor2_1 _08160_ (.A(_02587_),
    .B(_02560_),
    .Y(_00356_));
 sky130_fd_sc_hs__nor2_1 _08161_ (.A(_02585_),
    .B(_02584_),
    .Y(_02588_));
 sky130_fd_sc_hs__xnor2_1 _08162_ (.A(\u_fft.sched[54] ),
    .B(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hs__nor2_1 _08163_ (.A(_02589_),
    .B(_02560_),
    .Y(_00357_));
 sky130_fd_sc_hs__inv_2 _08164_ (.A(net2991),
    .Y(_02590_));
 sky130_fd_sc_hs__nor3_1 _08165_ (.A(net3780),
    .B(_00184_),
    .C(_02590_),
    .Y(_02591_));
 sky130_fd_sc_hs__o2bb2ai_1 _08166_ (.A1_N(net2960),
    .A2_N(_02591_),
    .B1(_00182_),
    .B2(_02560_),
    .Y(_00358_));
 sky130_fd_sc_hs__buf_2 place2133 (.A(_05473_),
    .X(net2133));
 sky130_fd_sc_hs__nand2_1 _08168_ (.A(_02559_),
    .B(\u_fft.sched[56] ),
    .Y(_02593_));
 sky130_fd_sc_hs__nand3_1 _08169_ (.A(net2960),
    .B(_00028_),
    .C(net2991),
    .Y(_02594_));
 sky130_fd_sc_hs__a21oi_1 _08170_ (.A1(_02593_),
    .A2(_02594_),
    .B1(net3780),
    .Y(_00359_));
 sky130_fd_sc_hs__xnor2_1 _08171_ (.A(_00027_),
    .B(_00188_),
    .Y(_02595_));
 sky130_fd_sc_hs__nor3_1 _08172_ (.A(_02590_),
    .B(_02595_),
    .C(_02559_),
    .Y(_02596_));
 sky130_fd_sc_hs__a21oi_1 _08173_ (.A1(\u_fft.sched[57] ),
    .A2(_02559_),
    .B1(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hs__nor2_1 _08174_ (.A(net3780),
    .B(_02597_),
    .Y(_00360_));
 sky130_fd_sc_hs__a21oi_1 _08175_ (.A1(_00188_),
    .A2(_00185_),
    .B1(_00187_),
    .Y(_02598_));
 sky130_fd_sc_hs__nand3_1 _08176_ (.A(_00026_),
    .B(_00186_),
    .C(_00188_),
    .Y(_02599_));
 sky130_fd_sc_hs__nand2_1 _08177_ (.A(_02598_),
    .B(_02599_),
    .Y(_02600_));
 sky130_fd_sc_hs__nand2_1 _08178_ (.A(_02600_),
    .B(_00190_),
    .Y(_02601_));
 sky130_fd_sc_hs__or2_1 _08179_ (.A(_00190_),
    .B(_02600_),
    .X(_02602_));
 sky130_fd_sc_hs__nand4_1 _08180_ (.A(net2960),
    .B(net2991),
    .C(_02601_),
    .D(_02602_),
    .Y(_02603_));
 sky130_fd_sc_hs__nand2_1 _08181_ (.A(_02559_),
    .B(\u_fft.sched[58] ),
    .Y(_02604_));
 sky130_fd_sc_hs__a21oi_1 _08182_ (.A1(_02603_),
    .A2(_02604_),
    .B1(net3780),
    .Y(_00361_));
 sky130_fd_sc_hs__a21oi_1 _08183_ (.A1(_00190_),
    .A2(_00187_),
    .B1(_00189_),
    .Y(_02605_));
 sky130_fd_sc_hs__nand3_1 _08184_ (.A(_00027_),
    .B(_00188_),
    .C(_00190_),
    .Y(_02606_));
 sky130_fd_sc_hs__nand2_1 _08185_ (.A(_02605_),
    .B(_02606_),
    .Y(_02607_));
 sky130_fd_sc_hs__xnor2_1 _08186_ (.A(_00192_),
    .B(_02607_),
    .Y(_02608_));
 sky130_fd_sc_hs__nor3_1 _08187_ (.A(_02590_),
    .B(_02608_),
    .C(_02559_),
    .Y(_02609_));
 sky130_fd_sc_hs__a21oi_1 _08188_ (.A1(\u_fft.sched[59] ),
    .A2(_02559_),
    .B1(_02609_),
    .Y(_02610_));
 sky130_fd_sc_hs__nor2_1 _08189_ (.A(net3780),
    .B(_02610_),
    .Y(_00362_));
 sky130_fd_sc_hs__inv_1 _08190_ (.A(_00194_),
    .Y(_02611_));
 sky130_fd_sc_hs__a21oi_1 _08191_ (.A1(_02600_),
    .A2(_00190_),
    .B1(_00189_),
    .Y(_02612_));
 sky130_fd_sc_hs__inv_1 _08192_ (.A(_02612_),
    .Y(_02613_));
 sky130_fd_sc_hs__a21oi_1 _08193_ (.A1(_02613_),
    .A2(_00192_),
    .B1(_00191_),
    .Y(_02614_));
 sky130_fd_sc_hs__nor2_1 _08194_ (.A(_02611_),
    .B(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hs__and2_1 _08195_ (.A(_02614_),
    .B(_02611_),
    .X(_02616_));
 sky130_fd_sc_hs__or4_1 _08196_ (.A(_02590_),
    .B(_02615_),
    .C(_02616_),
    .D(_02559_),
    .X(_02617_));
 sky130_fd_sc_hs__nand2_1 _08197_ (.A(_02559_),
    .B(\u_fft.sched[60] ),
    .Y(_02618_));
 sky130_fd_sc_hs__a21oi_1 _08198_ (.A1(_02617_),
    .A2(_02618_),
    .B1(net3780),
    .Y(_00363_));
 sky130_fd_sc_hs__a21oi_1 _08199_ (.A1(_02607_),
    .A2(_00192_),
    .B1(_00191_),
    .Y(_02619_));
 sky130_fd_sc_hs__o21bai_1 _08200_ (.A1(_02611_),
    .A2(_02619_),
    .B1_N(_00193_),
    .Y(_02620_));
 sky130_fd_sc_hs__nor2_1 _08201_ (.A(_00196_),
    .B(_02620_),
    .Y(_02621_));
 sky130_fd_sc_hs__nand2_1 _08202_ (.A(_02620_),
    .B(_00196_),
    .Y(_02622_));
 sky130_fd_sc_hs__nand3b_1 _08203_ (.A_N(_02621_),
    .B(net2991),
    .C(_02622_),
    .Y(_02623_));
 sky130_fd_sc_hs__nor2_1 _08204_ (.A(\u_fft.sched[61] ),
    .B(net2960),
    .Y(_02624_));
 sky130_fd_sc_hs__a211oi_1 _08205_ (.A1(net2960),
    .A2(_02623_),
    .B1(net3780),
    .C1(_02624_),
    .Y(_00364_));
 sky130_fd_sc_hs__nor2_1 _08206_ (.A(_00193_),
    .B(_02615_),
    .Y(_02625_));
 sky130_fd_sc_hs__inv_1 _08207_ (.A(_02625_),
    .Y(_02626_));
 sky130_fd_sc_hs__a21oi_1 _08208_ (.A1(_02626_),
    .A2(_00196_),
    .B1(_00195_),
    .Y(_02627_));
 sky130_fd_sc_hs__inv_1 _08209_ (.A(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hs__nor2_1 _08210_ (.A(_00198_),
    .B(_02628_),
    .Y(_02629_));
 sky130_fd_sc_hs__and2_1 _08211_ (.A(_02628_),
    .B(_00198_),
    .X(_02630_));
 sky130_fd_sc_hs__nor3_1 _08212_ (.A(_02629_),
    .B(_02630_),
    .C(_02590_),
    .Y(_02631_));
 sky130_fd_sc_hs__nand2_1 _08213_ (.A(_02631_),
    .B(net2960),
    .Y(_02632_));
 sky130_fd_sc_hs__nand2_1 _08214_ (.A(_02559_),
    .B(\u_fft.sched[62] ),
    .Y(_02633_));
 sky130_fd_sc_hs__a21oi_1 _08215_ (.A1(_02632_),
    .A2(_02633_),
    .B1(net3780),
    .Y(_00365_));
 sky130_fd_sc_hs__clkinv_1 _08216_ (.A(_00200_),
    .Y(_02634_));
 sky130_fd_sc_hs__nand2b_1 _08217_ (.A_N(_00195_),
    .B(_02622_),
    .Y(_02635_));
 sky130_fd_sc_hs__a21oi_1 _08218_ (.A1(_02635_),
    .A2(_00198_),
    .B1(_00197_),
    .Y(_02636_));
 sky130_fd_sc_hs__xnor2_1 _08219_ (.A(_02634_),
    .B(_02636_),
    .Y(_02637_));
 sky130_fd_sc_hs__nor3_1 _08220_ (.A(_02590_),
    .B(_02637_),
    .C(_02559_),
    .Y(_02638_));
 sky130_fd_sc_hs__a21oi_1 _08221_ (.A1(\u_fft.sched[63] ),
    .A2(_02559_),
    .B1(_02638_),
    .Y(_02639_));
 sky130_fd_sc_hs__nor2_1 _08222_ (.A(net3780),
    .B(_02639_),
    .Y(_00366_));
 sky130_fd_sc_hs__xnor2_1 _08223_ (.A(\u_fft.sched[39] ),
    .B(\u_fft.sched[64] ),
    .Y(_02640_));
 sky130_fd_sc_hs__nor2_1 _08224_ (.A(_00197_),
    .B(_02630_),
    .Y(_02641_));
 sky130_fd_sc_hs__o21bai_1 _08225_ (.A1(_02634_),
    .A2(_02641_),
    .B1_N(_00199_),
    .Y(_02642_));
 sky130_fd_sc_hs__xnor2_1 _08226_ (.A(_02640_),
    .B(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hs__nand3_1 _08227_ (.A(_02643_),
    .B(net2991),
    .C(net2960),
    .Y(_02644_));
 sky130_fd_sc_hs__nand2_1 _08228_ (.A(_02559_),
    .B(\u_fft.sched[64] ),
    .Y(_02645_));
 sky130_fd_sc_hs__a21oi_1 _08229_ (.A1(_02644_),
    .A2(_02645_),
    .B1(net3780),
    .Y(_00367_));
 sky130_fd_sc_hs__nor2_1 _08230_ (.A(\u_hamming_window.calc_pointer[0] ),
    .B(net3675),
    .Y(_00368_));
 sky130_fd_sc_hs__clkinv_1 _08231_ (.A(\u_hamming_window.calc_pointer[7] ),
    .Y(_02646_));
 sky130_fd_sc_hs__clkinv_1 _08232_ (.A(\u_hamming_window.calc_pointer[6] ),
    .Y(_02647_));
 sky130_fd_sc_hs__and2_1 _08233_ (.A(\u_hamming_window.calc_pointer[2] ),
    .B(_00239_),
    .X(_02648_));
 sky130_fd_sc_hs__nand3_1 _08234_ (.A(_02648_),
    .B(\u_hamming_window.calc_pointer[3] ),
    .C(\u_hamming_window.calc_pointer[4] ),
    .Y(_02649_));
 sky130_fd_sc_hs__nor2_1 _08235_ (.A(_05835_),
    .B(_02649_),
    .Y(_02650_));
 sky130_fd_sc_hs__inv_1 _08236_ (.A(_02650_),
    .Y(_02651_));
 sky130_fd_sc_hs__nor2_1 _08237_ (.A(_02647_),
    .B(_02651_),
    .Y(_02652_));
 sky130_fd_sc_hs__inv_1 _08238_ (.A(_02652_),
    .Y(_02653_));
 sky130_fd_sc_hs__nor2_1 _08239_ (.A(_02646_),
    .B(_02653_),
    .Y(_02654_));
 sky130_fd_sc_hs__inv_1 _08240_ (.A(\u_hamming_window.calc_pointer[9] ),
    .Y(_02655_));
 sky130_fd_sc_hs__inv_2 _08241_ (.A(\u_hamming_window.calc_pointer[8] ),
    .Y(_02656_));
 sky130_fd_sc_hs__nor2_1 _08242_ (.A(_02655_),
    .B(_02656_),
    .Y(_02657_));
 sky130_fd_sc_hs__a21oi_1 _08243_ (.A1(_02654_),
    .A2(_02657_),
    .B1(\u_hamming_window.calc_pointer[10] ),
    .Y(_02658_));
 sky130_fd_sc_hs__clkinv_1 _08244_ (.A(\u_hamming_window.calc_pointer[10] ),
    .Y(_02659_));
 sky130_fd_sc_hs__inv_1 _08245_ (.A(_02657_),
    .Y(_02660_));
 sky130_fd_sc_hs__inv_2 _08246_ (.A(_02654_),
    .Y(_02661_));
 sky130_fd_sc_hs__nor3_1 _08247_ (.A(_02659_),
    .B(_02660_),
    .C(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hs__nor3_1 _08248_ (.A(net3675),
    .B(_02658_),
    .C(_02662_),
    .Y(_00369_));
 sky130_fd_sc_hs__nor2_1 _08249_ (.A(_02646_),
    .B(_02656_),
    .Y(_02663_));
 sky130_fd_sc_hs__inv_2 _08250_ (.A(_02663_),
    .Y(_02664_));
 sky130_fd_sc_hs__clkinv_1 _08251_ (.A(\u_hamming_window.calc_pointer[4] ),
    .Y(_02665_));
 sky130_fd_sc_hs__nor3_1 _08252_ (.A(_05834_),
    .B(_00236_),
    .C(_00235_),
    .Y(_02666_));
 sky130_fd_sc_hs__nand2_1 _08253_ (.A(_02666_),
    .B(\u_hamming_window.calc_pointer[3] ),
    .Y(_02667_));
 sky130_fd_sc_hs__nor2_1 _08254_ (.A(_02665_),
    .B(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hs__nand2_1 _08255_ (.A(_02668_),
    .B(\u_hamming_window.calc_pointer[5] ),
    .Y(_02669_));
 sky130_fd_sc_hs__nor2_1 _08256_ (.A(_02647_),
    .B(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hs__inv_2 _08257_ (.A(_02670_),
    .Y(_02671_));
 sky130_fd_sc_hs__nor2_1 _08258_ (.A(_02664_),
    .B(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hs__inv_1 _08259_ (.A(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hs__nor2_1 _08260_ (.A(_02655_),
    .B(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hs__inv_1 _08261_ (.A(_02674_),
    .Y(_02675_));
 sky130_fd_sc_hs__clkinv_1 _08262_ (.A(\u_hamming_window.calc_pointer[11] ),
    .Y(_02676_));
 sky130_fd_sc_hs__nor2_1 _08263_ (.A(_02676_),
    .B(_02659_),
    .Y(_02677_));
 sky130_fd_sc_hs__inv_1 _08264_ (.A(_02677_),
    .Y(_02678_));
 sky130_fd_sc_hs__nor2_1 _08265_ (.A(_02678_),
    .B(_02675_),
    .Y(_02679_));
 sky130_fd_sc_hs__a2111oi_1 _08266_ (.A1(_02675_),
    .A2(_02676_),
    .B1(net3675),
    .C1(_05836_),
    .D1(_02679_),
    .Y(_00370_));
 sky130_fd_sc_hs__inv_1 _08267_ (.A(\u_hamming_window.calc_pointer[12] ),
    .Y(_02680_));
 sky130_fd_sc_hs__nand2_1 _08268_ (.A(_02662_),
    .B(\u_hamming_window.calc_pointer[11] ),
    .Y(_02681_));
 sky130_fd_sc_hs__buf_1 place2132 (.A(_05510_),
    .X(net2132));
 sky130_fd_sc_hs__o21ai_1 _08270_ (.A1(_02680_),
    .A2(_02681_),
    .B1(net3779),
    .Y(_02683_));
 sky130_fd_sc_hs__a21oi_1 _08271_ (.A1(_02680_),
    .A2(_02681_),
    .B1(_02683_),
    .Y(_00371_));
 sky130_fd_sc_hs__a21oi_1 _08272_ (.A1(_02679_),
    .A2(\u_hamming_window.calc_pointer[12] ),
    .B1(\u_hamming_window.calc_pointer[13] ),
    .Y(_02684_));
 sky130_fd_sc_hs__nand3_1 _08273_ (.A(_02679_),
    .B(\u_hamming_window.calc_pointer[13] ),
    .C(\u_hamming_window.calc_pointer[12] ),
    .Y(_02685_));
 sky130_fd_sc_hs__clkinv_1 _08274_ (.A(_02685_),
    .Y(_02686_));
 sky130_fd_sc_hs__nor3_1 _08275_ (.A(net3675),
    .B(_02684_),
    .C(_02686_),
    .Y(_00372_));
 sky130_fd_sc_hs__nor3_1 _08276_ (.A(_05828_),
    .B(_02680_),
    .C(_02681_),
    .Y(_02687_));
 sky130_fd_sc_hs__buf_1 place2131 (.A(_01732_),
    .X(net2131));
 sky130_fd_sc_hs__a21oi_1 _08278_ (.A1(_02687_),
    .A2(\u_hamming_window.calc_pointer[14] ),
    .B1(net3675),
    .Y(_02689_));
 sky130_fd_sc_hs__o21a_1 _08279_ (.A1(\u_hamming_window.calc_pointer[14] ),
    .A2(_02687_),
    .B1(_02689_),
    .X(_00373_));
 sky130_fd_sc_hs__nor2_1 _08280_ (.A(_05830_),
    .B(_05831_),
    .Y(_02690_));
 sky130_fd_sc_hs__inv_2 _08281_ (.A(_02690_),
    .Y(_02691_));
 sky130_fd_sc_hs__nor2_1 _08282_ (.A(_02691_),
    .B(_02685_),
    .Y(_02692_));
 sky130_fd_sc_hs__inv_1 _08283_ (.A(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hs__o2111a_1 _08284_ (.A1(\u_hamming_window.calc_pointer[15] ),
    .A2(_02686_),
    .B1(net3779),
    .C1(_05832_),
    .D1(_02693_),
    .X(_00374_));
 sky130_fd_sc_hs__clkinv_1 _08285_ (.A(\u_hamming_window.calc_pointer[16] ),
    .Y(_02694_));
 sky130_fd_sc_hs__nor3_1 _08286_ (.A(_05828_),
    .B(_02680_),
    .C(_02691_),
    .Y(_02695_));
 sky130_fd_sc_hs__nand4_1 _08287_ (.A(_02654_),
    .B(_02657_),
    .C(_02677_),
    .D(_02695_),
    .Y(_02696_));
 sky130_fd_sc_hs__nor2_1 _08288_ (.A(_02694_),
    .B(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hs__and2_1 _08289_ (.A(_02696_),
    .B(_02694_),
    .X(_02698_));
 sky130_fd_sc_hs__nor3_1 _08290_ (.A(_00589_),
    .B(_02697_),
    .C(_02698_),
    .Y(_00375_));
 sky130_fd_sc_hs__nor2_1 _08291_ (.A(_02694_),
    .B(_02693_),
    .Y(_02699_));
 sky130_fd_sc_hs__nor2_1 _08292_ (.A(\u_hamming_window.calc_pointer[17] ),
    .B(_02699_),
    .Y(_02700_));
 sky130_fd_sc_hs__nand2_1 _08293_ (.A(_02699_),
    .B(\u_hamming_window.calc_pointer[17] ),
    .Y(_02701_));
 sky130_fd_sc_hs__inv_2 _08294_ (.A(_02701_),
    .Y(_02702_));
 sky130_fd_sc_hs__nor3_1 _08295_ (.A(_00589_),
    .B(_02700_),
    .C(_02702_),
    .Y(_00376_));
 sky130_fd_sc_hs__clkinv_1 _08296_ (.A(\u_hamming_window.calc_pointer[18] ),
    .Y(_02703_));
 sky130_fd_sc_hs__nand2_1 _08297_ (.A(_02697_),
    .B(\u_hamming_window.calc_pointer[17] ),
    .Y(_02704_));
 sky130_fd_sc_hs__nor2_1 _08298_ (.A(_02703_),
    .B(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hs__inv_1 _08299_ (.A(_02705_),
    .Y(_02706_));
 sky130_fd_sc_hs__nand2_1 _08300_ (.A(_02706_),
    .B(net3779),
    .Y(_02707_));
 sky130_fd_sc_hs__a21oi_1 _08301_ (.A1(_02703_),
    .A2(_02704_),
    .B1(_02707_),
    .Y(_00377_));
 sky130_fd_sc_hs__clkinv_1 _08302_ (.A(\u_hamming_window.calc_pointer[19] ),
    .Y(_02708_));
 sky130_fd_sc_hs__nor2_1 _08303_ (.A(_02708_),
    .B(_02703_),
    .Y(_02709_));
 sky130_fd_sc_hs__nand2_1 _08304_ (.A(_02702_),
    .B(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hs__o2111a_1 _08305_ (.A1(\u_hamming_window.calc_pointer[19] ),
    .A2(_02702_),
    .B1(net3779),
    .C1(_05850_),
    .D1(_02710_),
    .X(_00378_));
 sky130_fd_sc_hs__and2_1 _08306_ (.A(net3779),
    .B(_00238_),
    .X(_00379_));
 sky130_fd_sc_hs__nor2_1 _08307_ (.A(_02708_),
    .B(_02706_),
    .Y(_02711_));
 sky130_fd_sc_hs__nor2_1 _08308_ (.A(\u_hamming_window.calc_pointer[20] ),
    .B(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hs__inv_1 _08309_ (.A(_02711_),
    .Y(_02713_));
 sky130_fd_sc_hs__nor2_1 _08310_ (.A(_00558_),
    .B(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hs__nor3_1 _08311_ (.A(_00589_),
    .B(_02712_),
    .C(_02714_),
    .Y(_00380_));
 sky130_fd_sc_hs__nor2_1 _08312_ (.A(_00558_),
    .B(_02710_),
    .Y(_02715_));
 sky130_fd_sc_hs__nor2_1 _08313_ (.A(\u_hamming_window.calc_pointer[21] ),
    .B(_02715_),
    .Y(_02716_));
 sky130_fd_sc_hs__nand2_1 _08314_ (.A(_02715_),
    .B(\u_hamming_window.calc_pointer[21] ),
    .Y(_02717_));
 sky130_fd_sc_hs__nor3b_1 _08315_ (.A(_00589_),
    .B(_02716_),
    .C_N(_02717_),
    .Y(_00381_));
 sky130_fd_sc_hs__nand2_1 _08316_ (.A(_02714_),
    .B(\u_hamming_window.calc_pointer[21] ),
    .Y(_02718_));
 sky130_fd_sc_hs__o21ai_1 _08317_ (.A1(_00560_),
    .A2(_02718_),
    .B1(net3779),
    .Y(_02719_));
 sky130_fd_sc_hs__a21oi_1 _08318_ (.A1(_00560_),
    .A2(_02718_),
    .B1(_02719_),
    .Y(_00382_));
 sky130_fd_sc_hs__nor2_1 _08319_ (.A(_00560_),
    .B(_02717_),
    .Y(_02720_));
 sky130_fd_sc_hs__inv_1 _08320_ (.A(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hs__o21ai_1 _08321_ (.A1(_00559_),
    .A2(_02721_),
    .B1(net3779),
    .Y(_02722_));
 sky130_fd_sc_hs__a21oi_1 _08322_ (.A1(_00559_),
    .A2(_02721_),
    .B1(_02722_),
    .Y(_00383_));
 sky130_fd_sc_hs__nand4_1 _08323_ (.A(_02714_),
    .B(\u_hamming_window.calc_pointer[21] ),
    .C(\u_hamming_window.calc_pointer[23] ),
    .D(\u_hamming_window.calc_pointer[22] ),
    .Y(_02723_));
 sky130_fd_sc_hs__o21ai_1 _08324_ (.A1(_05843_),
    .A2(_02723_),
    .B1(net3779),
    .Y(_02724_));
 sky130_fd_sc_hs__a21oi_1 _08325_ (.A1(_05843_),
    .A2(_02723_),
    .B1(_02724_),
    .Y(_00384_));
 sky130_fd_sc_hs__nor2_1 _08326_ (.A(_00559_),
    .B(_05843_),
    .Y(_02725_));
 sky130_fd_sc_hs__inv_1 _08327_ (.A(_02725_),
    .Y(_02726_));
 sky130_fd_sc_hs__nor2_1 _08328_ (.A(_00561_),
    .B(_02726_),
    .Y(_02727_));
 sky130_fd_sc_hs__a21oi_1 _08329_ (.A1(_02720_),
    .A2(_02725_),
    .B1(\u_hamming_window.calc_pointer[25] ),
    .Y(_02728_));
 sky130_fd_sc_hs__a211oi_1 _08330_ (.A1(_02720_),
    .A2(_02727_),
    .B1(_00589_),
    .C1(_02728_),
    .Y(_00385_));
 sky130_fd_sc_hs__nand2_1 _08331_ (.A(_02727_),
    .B(\u_hamming_window.calc_pointer[22] ),
    .Y(_02729_));
 sky130_fd_sc_hs__nor2_1 _08332_ (.A(_02729_),
    .B(_02718_),
    .Y(_02730_));
 sky130_fd_sc_hs__a21oi_1 _08333_ (.A1(_02730_),
    .A2(\u_hamming_window.calc_pointer[26] ),
    .B1(_00589_),
    .Y(_02731_));
 sky130_fd_sc_hs__o21a_1 _08334_ (.A1(\u_hamming_window.calc_pointer[26] ),
    .A2(_02730_),
    .B1(_02731_),
    .X(_00386_));
 sky130_fd_sc_hs__nand4_1 _08335_ (.A(_02720_),
    .B(\u_hamming_window.calc_pointer[25] ),
    .C(\u_hamming_window.calc_pointer[26] ),
    .D(_02725_),
    .Y(_02732_));
 sky130_fd_sc_hs__nor2_1 _08336_ (.A(_05840_),
    .B(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hs__inv_1 _08337_ (.A(_02733_),
    .Y(_02734_));
 sky130_fd_sc_hs__nand2_1 _08338_ (.A(_02734_),
    .B(net3779),
    .Y(_02735_));
 sky130_fd_sc_hs__a21oi_1 _08339_ (.A1(_05840_),
    .A2(_02732_),
    .B1(_02735_),
    .Y(_00387_));
 sky130_fd_sc_hs__nor2_1 _08340_ (.A(_05839_),
    .B(_00558_),
    .Y(_02736_));
 sky130_fd_sc_hs__nor2_1 _08341_ (.A(_05840_),
    .B(_05841_),
    .Y(_02737_));
 sky130_fd_sc_hs__nand4_1 _08342_ (.A(_02727_),
    .B(\u_hamming_window.calc_pointer[22] ),
    .C(_02736_),
    .D(_02737_),
    .Y(_02738_));
 sky130_fd_sc_hs__nor3_1 _08343_ (.A(_05845_),
    .B(_02738_),
    .C(_02713_),
    .Y(_02739_));
 sky130_fd_sc_hs__o21a_1 _08344_ (.A1(_02738_),
    .A2(_02713_),
    .B1(_05845_),
    .X(_02740_));
 sky130_fd_sc_hs__nor3_1 _08345_ (.A(_00589_),
    .B(_02739_),
    .C(_02740_),
    .Y(_00388_));
 sky130_fd_sc_hs__nor2_1 _08346_ (.A(_05845_),
    .B(_02734_),
    .Y(_02741_));
 sky130_fd_sc_hs__nor2_1 _08347_ (.A(\u_hamming_window.calc_pointer[29] ),
    .B(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hs__nand2_1 _08348_ (.A(_02741_),
    .B(\u_hamming_window.calc_pointer[29] ),
    .Y(_02743_));
 sky130_fd_sc_hs__clkinv_1 _08349_ (.A(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hs__nor3_1 _08350_ (.A(_00589_),
    .B(_02742_),
    .C(_02744_),
    .Y(_00389_));
 sky130_fd_sc_hs__nor2_1 _08351_ (.A(\u_hamming_window.calc_pointer[2] ),
    .B(_00239_),
    .Y(_02745_));
 sky130_fd_sc_hs__nor3_1 _08352_ (.A(net3675),
    .B(_02745_),
    .C(_02648_),
    .Y(_00390_));
 sky130_fd_sc_hs__nand3_1 _08353_ (.A(_02730_),
    .B(\u_hamming_window.calc_pointer[26] ),
    .C(\u_hamming_window.calc_pointer[29] ),
    .Y(_02746_));
 sky130_fd_sc_hs__nor3_1 _08354_ (.A(_05840_),
    .B(_05845_),
    .C(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hs__xnor2_1 _08355_ (.A(\u_hamming_window.calc_pointer[30] ),
    .B(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hs__nor2_1 _08356_ (.A(net3675),
    .B(_02748_),
    .Y(_00391_));
 sky130_fd_sc_hs__nor3b_1 _08357_ (.A(_05846_),
    .B(_02743_),
    .C_N(\u_hamming_window.calc_pointer[31] ),
    .Y(_02749_));
 sky130_fd_sc_hs__a21oi_1 _08358_ (.A1(_02744_),
    .A2(\u_hamming_window.calc_pointer[30] ),
    .B1(\u_hamming_window.calc_pointer[31] ),
    .Y(_02750_));
 sky130_fd_sc_hs__nor3_1 _08359_ (.A(_00589_),
    .B(_02749_),
    .C(_02750_),
    .Y(_00392_));
 sky130_fd_sc_hs__nor2_1 _08360_ (.A(\u_hamming_window.calc_pointer[3] ),
    .B(_02666_),
    .Y(_02751_));
 sky130_fd_sc_hs__nor3b_1 _08361_ (.A(net3675),
    .B(_02751_),
    .C_N(_02667_),
    .Y(_00393_));
 sky130_fd_sc_hs__a21oi_1 _08362_ (.A1(_02648_),
    .A2(\u_hamming_window.calc_pointer[3] ),
    .B1(\u_hamming_window.calc_pointer[4] ),
    .Y(_02752_));
 sky130_fd_sc_hs__nor3b_1 _08363_ (.A(net3675),
    .B(_02752_),
    .C_N(_02649_),
    .Y(_00394_));
 sky130_fd_sc_hs__nor2_1 _08364_ (.A(\u_hamming_window.calc_pointer[5] ),
    .B(_02668_),
    .Y(_02753_));
 sky130_fd_sc_hs__nor3b_1 _08365_ (.A(net3675),
    .B(_02753_),
    .C_N(_02669_),
    .Y(_00395_));
 sky130_fd_sc_hs__nor2_1 _08366_ (.A(\u_hamming_window.calc_pointer[6] ),
    .B(_02650_),
    .Y(_02754_));
 sky130_fd_sc_hs__nor3_1 _08367_ (.A(net3675),
    .B(_02754_),
    .C(_02652_),
    .Y(_00396_));
 sky130_fd_sc_hs__o21ai_1 _08368_ (.A1(_02646_),
    .A2(_02671_),
    .B1(net3779),
    .Y(_02755_));
 sky130_fd_sc_hs__a21oi_1 _08369_ (.A1(_02646_),
    .A2(_02671_),
    .B1(_02755_),
    .Y(_00397_));
 sky130_fd_sc_hs__o21ai_1 _08370_ (.A1(_02656_),
    .A2(_02661_),
    .B1(net3779),
    .Y(_02756_));
 sky130_fd_sc_hs__a21oi_1 _08371_ (.A1(_02656_),
    .A2(_02661_),
    .B1(_02756_),
    .Y(_00398_));
 sky130_fd_sc_hs__nor2_1 _08372_ (.A(\u_hamming_window.calc_pointer[9] ),
    .B(_02672_),
    .Y(_02757_));
 sky130_fd_sc_hs__nor3_1 _08373_ (.A(net3675),
    .B(_02757_),
    .C(_02674_),
    .Y(_00399_));
 sky130_fd_sc_hs__nor2_1 _08374_ (.A(_05774_),
    .B(_00669_),
    .Y(_00400_));
 sky130_fd_sc_hs__nor2_1 _08375_ (.A(\u_hamming_window.hamming_state[2] ),
    .B(\u_hamming_window.hamming_state[1] ),
    .Y(_02758_));
 sky130_fd_sc_hs__nor2_1 _08376_ (.A(\u_hamming_window.hamming_state[0] ),
    .B(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hs__o22a_2 _08377_ (.A1(_00567_),
    .A2(_02759_),
    .B1(_02237_),
    .B2(_00588_),
    .X(_02760_));
 sky130_fd_sc_hs__and2_2 _08378_ (.A(net1844),
    .B(_02760_),
    .X(_02761_));
 sky130_fd_sc_hs__nor2_2 _08379_ (.A(\u_hamming_window.frame_ptr[0] ),
    .B(_02761_),
    .Y(_02762_));
 sky130_fd_sc_hs__bufbuf_8 place2130 (.A(net4932),
    .X(net2130));
 sky130_fd_sc_hs__nand3_1 _08381_ (.A(net1844),
    .B(\u_hamming_window.frame_ptr[0] ),
    .C(_02760_),
    .Y(_02764_));
 sky130_fd_sc_hs__a31oi_1 _08382_ (.A1(_02758_),
    .A2(\u_hamming_window.hamming_state[0] ),
    .A3(start_hamming),
    .B1(net3782),
    .Y(_02765_));
 sky130_fd_sc_hs__nand2_1 _08383_ (.A(_02764_),
    .B(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hs__nor2_1 _08384_ (.A(_02762_),
    .B(_02766_),
    .Y(_00401_));
 sky130_fd_sc_hs__nor2_2 _08385_ (.A(\u_hamming_window.frame_ptr[1] ),
    .B(_02761_),
    .Y(_02767_));
 sky130_fd_sc_hs__nand3b_1 _08386_ (.A_N(_00204_),
    .B(net1844),
    .C(_02760_),
    .Y(_02768_));
 sky130_fd_sc_hs__nand2_1 _08387_ (.A(_02768_),
    .B(_02765_),
    .Y(_02769_));
 sky130_fd_sc_hs__nor2_1 _08388_ (.A(_02767_),
    .B(_02769_),
    .Y(_00402_));
 sky130_fd_sc_hs__nand2_2 _08389_ (.A(net1844),
    .B(_02760_),
    .Y(_02770_));
 sky130_fd_sc_hs__nand2_2 _08390_ (.A(net1841),
    .B(\u_hamming_window.frame_ptr[2] ),
    .Y(_02771_));
 sky130_fd_sc_hs__xnor2_1 _08391_ (.A(\u_hamming_window.frame_ptr[2] ),
    .B(_00203_),
    .Y(_02772_));
 sky130_fd_sc_hs__nor2_1 _08392_ (.A(_02758_),
    .B(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hs__nand3_1 _08393_ (.A(net1844),
    .B(_02760_),
    .C(_02773_),
    .Y(_02774_));
 sky130_fd_sc_hs__a21boi_1 _08394_ (.A1(_02774_),
    .A2(_02771_),
    .B1_N(net211),
    .Y(_00403_));
 sky130_fd_sc_hs__nand2_2 _08395_ (.A(net1841),
    .B(\u_hamming_window.frame_ptr[3] ),
    .Y(_02775_));
 sky130_fd_sc_hs__nand3_1 _08396_ (.A(\u_hamming_window.frame_ptr[0] ),
    .B(\u_hamming_window.frame_ptr[2] ),
    .C(\u_hamming_window.frame_ptr[1] ),
    .Y(_02776_));
 sky130_fd_sc_hs__xor2_1 _08397_ (.A(\u_hamming_window.frame_ptr[3] ),
    .B(_02776_),
    .X(_02777_));
 sky130_fd_sc_hs__nor2_1 _08398_ (.A(_02758_),
    .B(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hs__nand3_1 _08399_ (.A(net1844),
    .B(_02760_),
    .C(_02778_),
    .Y(_02779_));
 sky130_fd_sc_hs__a21boi_2 _08400_ (.A1(_02779_),
    .A2(_02775_),
    .B1_N(net211),
    .Y(_00404_));
 sky130_fd_sc_hs__nand2_2 _08401_ (.A(net1841),
    .B(\u_hamming_window.frame_ptr[4] ),
    .Y(_02780_));
 sky130_fd_sc_hs__clkinv_1 _08402_ (.A(_00203_),
    .Y(_02781_));
 sky130_fd_sc_hs__nand2_1 _08403_ (.A(\u_hamming_window.frame_ptr[3] ),
    .B(\u_hamming_window.frame_ptr[2] ),
    .Y(_02782_));
 sky130_fd_sc_hs__nor2_1 _08404_ (.A(_02781_),
    .B(_02782_),
    .Y(_02783_));
 sky130_fd_sc_hs__xnor2_1 _08405_ (.A(\u_hamming_window.frame_ptr[4] ),
    .B(_02783_),
    .Y(_02784_));
 sky130_fd_sc_hs__nor2_1 _08406_ (.A(_02758_),
    .B(_02784_),
    .Y(_02785_));
 sky130_fd_sc_hs__nand3_1 _08407_ (.A(net5041),
    .B(_02760_),
    .C(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hs__a21boi_2 _08408_ (.A1(_02780_),
    .A2(_02786_),
    .B1_N(net211),
    .Y(_00405_));
 sky130_fd_sc_hs__nand3_1 _08409_ (.A(net5040),
    .B(_00587_),
    .C(_02760_),
    .Y(_02787_));
 sky130_fd_sc_hs__nand2_1 _08410_ (.A(_02787_),
    .B(_02765_),
    .Y(_02788_));
 sky130_fd_sc_hs__inv_1 _08411_ (.A(_00586_),
    .Y(_02789_));
 sky130_fd_sc_hs__nand3_2 _08412_ (.A(net5040),
    .B(_02789_),
    .C(_02760_),
    .Y(_02790_));
 sky130_fd_sc_hs__and2_2 _08413_ (.A(_00582_),
    .B(_02790_),
    .X(_02791_));
 sky130_fd_sc_hs__nor2_2 _08414_ (.A(_02791_),
    .B(_02788_),
    .Y(_00406_));
 sky130_fd_sc_hs__nand2_2 _08415_ (.A(net1841),
    .B(\u_hamming_window.frame_ptr[6] ),
    .Y(_02792_));
 sky130_fd_sc_hs__nor4_1 _08416_ (.A(_00582_),
    .B(_00583_),
    .C(_02781_),
    .D(_02782_),
    .Y(_02793_));
 sky130_fd_sc_hs__xnor2_1 _08417_ (.A(\u_hamming_window.frame_ptr[6] ),
    .B(_02793_),
    .Y(_02794_));
 sky130_fd_sc_hs__nor2_1 _08418_ (.A(_02758_),
    .B(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hs__nand3_1 _08419_ (.A(net5041),
    .B(_02760_),
    .C(_02795_),
    .Y(_02796_));
 sky130_fd_sc_hs__a21boi_2 _08420_ (.A1(_02796_),
    .A2(_02792_),
    .B1_N(net211),
    .Y(_00407_));
 sky130_fd_sc_hs__nand2_1 _08421_ (.A(net1841),
    .B(\u_hamming_window.frame_ptr[7] ),
    .Y(_02797_));
 sky130_fd_sc_hs__nand2_1 _08422_ (.A(_00587_),
    .B(\u_hamming_window.frame_ptr[6] ),
    .Y(_02798_));
 sky130_fd_sc_hs__xor2_1 _08423_ (.A(\u_hamming_window.frame_ptr[7] ),
    .B(_02798_),
    .X(_02799_));
 sky130_fd_sc_hs__nor2_1 _08424_ (.A(_02758_),
    .B(_02799_),
    .Y(_02800_));
 sky130_fd_sc_hs__nand3_1 _08425_ (.A(net5040),
    .B(_02760_),
    .C(_02800_),
    .Y(_02801_));
 sky130_fd_sc_hs__a21boi_1 _08426_ (.A1(_02797_),
    .A2(_02801_),
    .B1_N(net211),
    .Y(_00408_));
 sky130_fd_sc_hs__nand2_1 _08427_ (.A(net1841),
    .B(\u_hamming_window.frame_ptr[8] ),
    .Y(_02802_));
 sky130_fd_sc_hs__nor3_1 _08428_ (.A(_00582_),
    .B(_00583_),
    .C(_00581_),
    .Y(_02803_));
 sky130_fd_sc_hs__nand2_1 _08429_ (.A(_02803_),
    .B(_02783_),
    .Y(_02804_));
 sky130_fd_sc_hs__xor2_1 _08430_ (.A(\u_hamming_window.frame_ptr[8] ),
    .B(_02804_),
    .X(_02805_));
 sky130_fd_sc_hs__nor2_1 _08431_ (.A(_02758_),
    .B(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hs__nand3_1 _08432_ (.A(net5041),
    .B(_02760_),
    .C(_02806_),
    .Y(_02807_));
 sky130_fd_sc_hs__a21boi_1 _08433_ (.A1(_02802_),
    .A2(_02807_),
    .B1_N(net211),
    .Y(_00409_));
 sky130_fd_sc_hs__nor2_1 _08434_ (.A(net3782),
    .B(_00568_),
    .Y(_00410_));
 sky130_fd_sc_hs__nand2_1 _08435_ (.A(_05816_),
    .B(\u_mel.state[1] ),
    .Y(_02808_));
 sky130_fd_sc_hs__o211ai_1 _08436_ (.A1(\u_mel.state[2] ),
    .A2(\u_mel.state[1] ),
    .B1(_05824_),
    .C1(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hs__o21ai_1 _08437_ (.A1(\u_mel.k_next[0] ),
    .A2(_02809_),
    .B1(net211),
    .Y(_02810_));
 sky130_fd_sc_hs__a21oi_1 _08438_ (.A1(\u_mel.k_next[0] ),
    .A2(_02809_),
    .B1(_02810_),
    .Y(_00411_));
 sky130_fd_sc_hs__o21ai_1 _08439_ (.A1(\u_mel.k_next[1] ),
    .A2(_02809_),
    .B1(net211),
    .Y(_02811_));
 sky130_fd_sc_hs__a21oi_1 _08440_ (.A1(_00240_),
    .A2(_02809_),
    .B1(_02811_),
    .Y(_00412_));
 sky130_fd_sc_hs__nor2b_1 _08441_ (.A(_02809_),
    .B_N(_00242_),
    .Y(_02812_));
 sky130_fd_sc_hs__nor2_1 _08442_ (.A(\u_mel.k[2] ),
    .B(_02812_),
    .Y(_02813_));
 sky130_fd_sc_hs__nand2_1 _08443_ (.A(_02812_),
    .B(\u_mel.k[2] ),
    .Y(_02814_));
 sky130_fd_sc_hs__nor3b_1 _08444_ (.A(net3781),
    .B(_02813_),
    .C_N(_02814_),
    .Y(_00413_));
 sky130_fd_sc_hs__nand2_1 _08445_ (.A(\u_mel.k[2] ),
    .B(\u_mel.k[1] ),
    .Y(_02815_));
 sky130_fd_sc_hs__nor3_1 _08446_ (.A(\u_mel.k_next[0] ),
    .B(_02815_),
    .C(_02809_),
    .Y(_02816_));
 sky130_fd_sc_hs__nor2_1 _08447_ (.A(\u_mel.k[3] ),
    .B(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hs__nand2_1 _08448_ (.A(_02816_),
    .B(\u_mel.k[3] ),
    .Y(_02818_));
 sky130_fd_sc_hs__nor3b_1 _08449_ (.A(net3781),
    .B(_02817_),
    .C_N(_02818_),
    .Y(_00414_));
 sky130_fd_sc_hs__and3_1 _08450_ (.A(_02812_),
    .B(\u_mel.k[3] ),
    .C(\u_mel.k[2] ),
    .X(_02819_));
 sky130_fd_sc_hs__nor2_1 _08451_ (.A(\u_mel.k[4] ),
    .B(_02819_),
    .Y(_02820_));
 sky130_fd_sc_hs__nand2_1 _08452_ (.A(_02819_),
    .B(\u_mel.k[4] ),
    .Y(_02821_));
 sky130_fd_sc_hs__nor3b_1 _08453_ (.A(net3781),
    .B(_02820_),
    .C_N(_02821_),
    .Y(_00415_));
 sky130_fd_sc_hs__nor2_1 _08454_ (.A(_05809_),
    .B(_02818_),
    .Y(_02822_));
 sky130_fd_sc_hs__nor2_1 _08455_ (.A(\u_mel.k[5] ),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hs__nand2_1 _08456_ (.A(_02822_),
    .B(\u_mel.k[5] ),
    .Y(_02824_));
 sky130_fd_sc_hs__clkinv_1 _08457_ (.A(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hs__nor3_1 _08458_ (.A(net3781),
    .B(_02823_),
    .C(_02825_),
    .Y(_00416_));
 sky130_fd_sc_hs__nor2_1 _08459_ (.A(_05808_),
    .B(_02821_),
    .Y(_02826_));
 sky130_fd_sc_hs__nor2_1 _08460_ (.A(\u_mel.k[6] ),
    .B(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hs__nand2_1 _08461_ (.A(_02826_),
    .B(\u_mel.k[6] ),
    .Y(_02828_));
 sky130_fd_sc_hs__nor3b_1 _08462_ (.A(net3781),
    .B(_02827_),
    .C_N(_02828_),
    .Y(_00417_));
 sky130_fd_sc_hs__nor3_1 _08463_ (.A(_05811_),
    .B(_05812_),
    .C(_02824_),
    .Y(_02829_));
 sky130_fd_sc_hs__a21oi_1 _08464_ (.A1(_02825_),
    .A2(\u_mel.k[6] ),
    .B1(\u_mel.k[7] ),
    .Y(_02830_));
 sky130_fd_sc_hs__nor3_1 _08465_ (.A(net3781),
    .B(_02829_),
    .C(_02830_),
    .Y(_00418_));
 sky130_fd_sc_hs__nor3_1 _08466_ (.A(_05811_),
    .B(_05813_),
    .C(_02828_),
    .Y(_02831_));
 sky130_fd_sc_hs__a31oi_1 _08467_ (.A1(_02826_),
    .A2(\u_mel.k[7] ),
    .A3(\u_mel.k[6] ),
    .B1(\u_mel.k[8] ),
    .Y(_02832_));
 sky130_fd_sc_hs__nor3_1 _08468_ (.A(net3781),
    .B(_02831_),
    .C(_02832_),
    .Y(_00419_));
 sky130_fd_sc_hs__nor2_1 _08469_ (.A(net3781),
    .B(_05819_),
    .Y(_00420_));
 sky130_fd_sc_hs__inv_2 _08470_ (.A(mel_valid),
    .Y(_02833_));
 sky130_fd_sc_hs__nor2_1 _08471_ (.A(\u_mel.state[0] ),
    .B(mel_valid),
    .Y(_02834_));
 sky130_fd_sc_hs__o21ai_1 _08472_ (.A1(_00205_),
    .A2(_02834_),
    .B1(net211),
    .Y(_02835_));
 sky130_fd_sc_hs__a21oi_1 _08473_ (.A1(_02833_),
    .A2(_00205_),
    .B1(_02835_),
    .Y(_00421_));
 sky130_fd_sc_hs__nand2_1 _08474_ (.A(_02834_),
    .B(\mel_ptr[1] ),
    .Y(_02836_));
 sky130_fd_sc_hs__nand2_1 _08475_ (.A(mel_valid),
    .B(_00208_),
    .Y(_02837_));
 sky130_fd_sc_hs__a21oi_1 _08476_ (.A1(_02836_),
    .A2(_02837_),
    .B1(net3781),
    .Y(_00422_));
 sky130_fd_sc_hs__nand2_1 _08477_ (.A(_02834_),
    .B(\mel_ptr[2] ),
    .Y(_02838_));
 sky130_fd_sc_hs__nand2_1 _08478_ (.A(\mel_ptr[2] ),
    .B(_00209_),
    .Y(_02839_));
 sky130_fd_sc_hs__nand2_1 _08479_ (.A(_02839_),
    .B(mel_valid),
    .Y(_02840_));
 sky130_fd_sc_hs__o21ai_1 _08480_ (.A1(\mel_ptr[2] ),
    .A2(_00209_),
    .B1(net211),
    .Y(_02841_));
 sky130_fd_sc_hs__a21oi_1 _08481_ (.A1(_02838_),
    .A2(_02840_),
    .B1(_02841_),
    .Y(_00423_));
 sky130_fd_sc_hs__nor4_1 _08482_ (.A(_05818_),
    .B(_02833_),
    .C(_00206_),
    .D(_00205_),
    .Y(_02842_));
 sky130_fd_sc_hs__nand2_1 _08483_ (.A(_02833_),
    .B(\u_mel.state[0] ),
    .Y(_02843_));
 sky130_fd_sc_hs__a21oi_1 _08484_ (.A1(\mel_ptr[3] ),
    .A2(_02843_),
    .B1(_02842_),
    .Y(_02844_));
 sky130_fd_sc_hs__a211oi_1 _08485_ (.A1(\mel_ptr[3] ),
    .A2(_02842_),
    .B1(net3781),
    .C1(_02844_),
    .Y(_00424_));
 sky130_fd_sc_hs__nor2_1 _08486_ (.A(_05801_),
    .B(_02839_),
    .Y(_02845_));
 sky130_fd_sc_hs__a22oi_1 _08487_ (.A1(_02843_),
    .A2(\mel_ptr[4] ),
    .B1(mel_valid),
    .B2(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hs__a311oi_1 _08488_ (.A1(\mel_ptr[4] ),
    .A2(mel_valid),
    .A3(_02845_),
    .B1(net3781),
    .C1(_02846_),
    .Y(_00425_));
 sky130_fd_sc_hs__nor3b_1 _08489_ (.A(_05801_),
    .B(_05802_),
    .C_N(_02842_),
    .Y(_02847_));
 sky130_fd_sc_hs__a21oi_1 _08490_ (.A1(\mel_ptr[5] ),
    .A2(_02843_),
    .B1(_02847_),
    .Y(_02848_));
 sky130_fd_sc_hs__a211oi_1 _08491_ (.A1(\mel_ptr[5] ),
    .A2(_02847_),
    .B1(net3781),
    .C1(_02848_),
    .Y(_00426_));
 sky130_fd_sc_hs__nand3_1 _08492_ (.A(_00648_),
    .B(_00225_),
    .C(_00640_),
    .Y(_02849_));
 sky130_fd_sc_hs__o311ai_1 _08493_ (.A1(_00638_),
    .A2(_00630_),
    .A3(_02849_),
    .B1(\u_window_buffer.current_state[2] ),
    .C1(_00612_),
    .Y(_02850_));
 sky130_fd_sc_hs__a21oi_1 _08494_ (.A1(_02850_),
    .A2(_00655_),
    .B1(net3782),
    .Y(_00427_));
 sky130_fd_sc_hs__nor2_1 _08495_ (.A(_02224_),
    .B(net3615),
    .Y(_02851_));
 sky130_fd_sc_hs__inv_2 _08496_ (.A(_02851_),
    .Y(_02852_));
 sky130_fd_sc_hs__nand2_1 _08497_ (.A(net3775),
    .B(net3776),
    .Y(_02853_));
 sky130_fd_sc_hs__inv_1 _08498_ (.A(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hs__nand2_1 _08499_ (.A(net3749),
    .B(net3748),
    .Y(_02855_));
 sky130_fd_sc_hs__nand2_1 _08500_ (.A(_02855_),
    .B(_02193_),
    .Y(_02856_));
 sky130_fd_sc_hs__nand3_2 _08501_ (.A(_02192_),
    .B(_02854_),
    .C(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hs__nor2_2 _08502_ (.A(_02188_),
    .B(_02857_),
    .Y(_02858_));
 sky130_fd_sc_hs__nand2_1 _08503_ (.A(_02214_),
    .B(_02198_),
    .Y(_02859_));
 sky130_fd_sc_hs__inv_2 _08504_ (.A(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hs__nand4_2 _08505_ (.A(_02858_),
    .B(net3766),
    .C(_02860_),
    .D(_02211_),
    .Y(_02861_));
 sky130_fd_sc_hs__nor2_2 _08506_ (.A(net3621),
    .B(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hs__nand3_1 _08507_ (.A(_02862_),
    .B(net3761),
    .C(_02202_),
    .Y(_02863_));
 sky130_fd_sc_hs__nor2_4 _08508_ (.A(net3612),
    .B(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hs__nand2_4 _08509_ (.A(_02864_),
    .B(net3759),
    .Y(_02865_));
 sky130_fd_sc_hs__nor3_2 _08510_ (.A(net3611),
    .B(_02852_),
    .C(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hs__nand2_1 _08511_ (.A(_02866_),
    .B(net3755),
    .Y(_02867_));
 sky130_fd_sc_hs__xor2_2 _08512_ (.A(net3753),
    .B(_02867_),
    .X(_02868_));
 sky130_fd_sc_hs__nand3_4 _08513_ (.A(net3336),
    .B(net3446),
    .C(net3301),
    .Y(_02869_));
 sky130_fd_sc_hs__or2_4 _08514_ (.A(_02207_),
    .B(_02869_),
    .X(_02870_));
 sky130_fd_sc_hs__or2_4 _08515_ (.A(_02203_),
    .B(_02870_),
    .X(_02871_));
 sky130_fd_sc_hs__nand3b_2 _08516_ (.A_N(_02871_),
    .B(net3760),
    .C(net3761),
    .Y(_02872_));
 sky130_fd_sc_hs__nor2_4 _08517_ (.A(_02872_),
    .B(net3614),
    .Y(_02873_));
 sky130_fd_sc_hs__nor2_1 _08518_ (.A(net3611),
    .B(net3385),
    .Y(_02874_));
 sky130_fd_sc_hs__nand2_1 _08519_ (.A(_02873_),
    .B(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hs__xor2_2 _08520_ (.A(net3755),
    .B(_02875_),
    .X(_02876_));
 sky130_fd_sc_hs__nand2_2 _08521_ (.A(_02873_),
    .B(net3758),
    .Y(_02877_));
 sky130_fd_sc_hs__xnor2_4 _08522_ (.A(_02877_),
    .B(net3610),
    .Y(_02878_));
 sky130_fd_sc_hs__nor2_1 _08523_ (.A(net3384),
    .B(net3130),
    .Y(_02879_));
 sky130_fd_sc_hs__o21bai_2 _08524_ (.A1(net3756),
    .A2(_02879_),
    .B1_N(net3085),
    .Y(_02880_));
 sky130_fd_sc_hs__xnor2_4 _08525_ (.A(net3615),
    .B(net3130),
    .Y(_02881_));
 sky130_fd_sc_hs__nand4_2 _08526_ (.A(net2988),
    .B(net5123),
    .C(_02880_),
    .D(net3084),
    .Y(_02882_));
 sky130_fd_sc_hs__xnor2_2 _08527_ (.A(net3614),
    .B(net3129),
    .Y(_02883_));
 sky130_fd_sc_hs__and2_1 _08528_ (.A(net3223),
    .B(net3613),
    .X(_02884_));
 sky130_fd_sc_hs__nor2_1 _08529_ (.A(net3179),
    .B(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hs__inv_1 _08530_ (.A(net3128),
    .Y(_02886_));
 sky130_fd_sc_hs__nand2_1 _08531_ (.A(net3082),
    .B(_02886_),
    .Y(_02887_));
 sky130_fd_sc_hs__xnor2_1 _08532_ (.A(net3766),
    .B(net3264),
    .Y(_02888_));
 sky130_fd_sc_hs__clkinv_1 _08533_ (.A(net3773),
    .Y(_02889_));
 sky130_fd_sc_hs__nor3_4 _08534_ (.A(_02889_),
    .B(_02188_),
    .C(net3383),
    .Y(_02890_));
 sky130_fd_sc_hs__nand3_2 _08535_ (.A(_02890_),
    .B(net3770),
    .C(net3771),
    .Y(_02891_));
 sky130_fd_sc_hs__nor3_4 _08536_ (.A(net3618),
    .B(net3617),
    .C(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hs__or2_1 _08537_ (.A(net3767),
    .B(_02892_),
    .X(_02893_));
 sky130_fd_sc_hs__nand2_1 _08538_ (.A(_02892_),
    .B(net3767),
    .Y(_02894_));
 sky130_fd_sc_hs__nand2_2 _08539_ (.A(_02893_),
    .B(_02894_),
    .Y(_02895_));
 sky130_fd_sc_hs__nand2_1 _08540_ (.A(net5176),
    .B(net3336),
    .Y(_02896_));
 sky130_fd_sc_hs__xnor2_1 _08541_ (.A(net3618),
    .B(_02896_),
    .Y(_02897_));
 sky130_fd_sc_hs__nand2_2 _08542_ (.A(_02895_),
    .B(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hs__xnor2_2 _08543_ (.A(net3616),
    .B(_02199_),
    .Y(_02899_));
 sky130_fd_sc_hs__xnor2_1 _08544_ (.A(net3771),
    .B(net3335),
    .Y(_02900_));
 sky130_fd_sc_hs__nand2_1 _08545_ (.A(_02899_),
    .B(net3297),
    .Y(_02901_));
 sky130_fd_sc_hs__xnor2_1 _08546_ (.A(net3628),
    .B(net3444),
    .Y(_02902_));
 sky130_fd_sc_hs__nor2_1 _08547_ (.A(net3751),
    .B(net3750),
    .Y(_02903_));
 sky130_fd_sc_hs__nand4_1 _08548_ (.A(_02903_),
    .B(_00210_),
    .C(_00211_),
    .D(net3749),
    .Y(_02904_));
 sky130_fd_sc_hs__nand2_1 _08549_ (.A(net3747),
    .B(net5183),
    .Y(_02905_));
 sky130_fd_sc_hs__and2_2 _08550_ (.A(net3389),
    .B(_02905_),
    .X(_02906_));
 sky130_fd_sc_hs__inv_2 _08551_ (.A(_02906_),
    .Y(_02907_));
 sky130_fd_sc_hs__nor3_2 _08552_ (.A(_00219_),
    .B(_02904_),
    .C(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hs__nand2b_1 _08553_ (.A_N(_02902_),
    .B(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hs__xnor2_1 _08554_ (.A(net3607),
    .B(net5195),
    .Y(_02910_));
 sky130_fd_sc_hs__clkinv_1 _08555_ (.A(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hs__a21oi_1 _08556_ (.A1(net3627),
    .A2(net3447),
    .B1(net3628),
    .Y(_02912_));
 sky130_fd_sc_hs__xnor2_1 _08557_ (.A(net3629),
    .B(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hs__inv_1 _08558_ (.A(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hs__nand3_1 _08559_ (.A(_02856_),
    .B(net3745),
    .C(net3746),
    .Y(_02915_));
 sky130_fd_sc_hs__xor2_1 _08560_ (.A(net3776),
    .B(_02915_),
    .X(_02916_));
 sky130_fd_sc_hs__nand2_2 _08561_ (.A(_02914_),
    .B(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hs__xnor2_2 _08562_ (.A(net3775),
    .B(net3337),
    .Y(_02918_));
 sky130_fd_sc_hs__inv_2 _08563_ (.A(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hs__xnor2_2 _08564_ (.A(net3630),
    .B(net3383),
    .Y(_02920_));
 sky130_fd_sc_hs__nand2_1 _08565_ (.A(_02919_),
    .B(_02920_),
    .Y(_02921_));
 sky130_fd_sc_hs__nor2_2 _08566_ (.A(_02917_),
    .B(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hs__nand3b_1 _08567_ (.A_N(_02909_),
    .B(_02922_),
    .C(_02911_),
    .Y(_02923_));
 sky130_fd_sc_hs__nor2_4 _08568_ (.A(_02923_),
    .B(_02901_),
    .Y(_02924_));
 sky130_fd_sc_hs__xnor2_2 _08569_ (.A(net3617),
    .B(net3298),
    .Y(_02925_));
 sky130_fd_sc_hs__nand2_1 _08570_ (.A(_02924_),
    .B(net3258),
    .Y(_02926_));
 sky130_fd_sc_hs__nor3_2 _08571_ (.A(_02888_),
    .B(_02898_),
    .C(_02926_),
    .Y(_02927_));
 sky130_fd_sc_hs__and2_1 _08572_ (.A(net3299),
    .B(net3621),
    .X(_02928_));
 sky130_fd_sc_hs__nor2_1 _08573_ (.A(net3265),
    .B(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hs__inv_1 _08574_ (.A(_02929_),
    .Y(_02930_));
 sky130_fd_sc_hs__xnor2_2 _08575_ (.A(net3761),
    .B(net3178),
    .Y(_02931_));
 sky130_fd_sc_hs__nor4_1 _08576_ (.A(net3622),
    .B(net3621),
    .C(net3620),
    .D(net3619),
    .Y(_02932_));
 sky130_fd_sc_hs__nand2_1 _08577_ (.A(net3263),
    .B(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hs__xnor2_2 _08578_ (.A(net3624),
    .B(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hs__xnor2_2 _08579_ (.A(net3623),
    .B(net3222),
    .Y(_02935_));
 sky130_fd_sc_hs__nand2_1 _08580_ (.A(_02934_),
    .B(_02935_),
    .Y(_02936_));
 sky130_fd_sc_hs__nor2_2 _08581_ (.A(_02931_),
    .B(_02936_),
    .Y(_02937_));
 sky130_fd_sc_hs__nand3_2 _08582_ (.A(net2985),
    .B(_02930_),
    .C(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hs__o21a_1 _08583_ (.A1(_02938_),
    .A2(_02887_),
    .B1(_02232_),
    .X(_02939_));
 sky130_fd_sc_hs__a21oi_4 _08584_ (.A1(_02882_),
    .A2(net3086),
    .B1(_02939_),
    .Y(_02940_));
 sky130_fd_sc_hs__xor2_4 _08585_ (.A(_02940_),
    .B(net2990),
    .X(_02941_));
 sky130_fd_sc_hs__nor2_2 _08586_ (.A(_02885_),
    .B(_02931_),
    .Y(_02942_));
 sky130_fd_sc_hs__nand3_1 _08587_ (.A(_02883_),
    .B(_02942_),
    .C(_02881_),
    .Y(_02943_));
 sky130_fd_sc_hs__nand2_2 _08588_ (.A(_02878_),
    .B(_02880_),
    .Y(_02944_));
 sky130_fd_sc_hs__nand2_1 _08589_ (.A(_02868_),
    .B(_02876_),
    .Y(_02945_));
 sky130_fd_sc_hs__nor3_4 _08590_ (.A(_02943_),
    .B(_02944_),
    .C(_02945_),
    .Y(_02946_));
 sky130_fd_sc_hs__nand2_2 _08591_ (.A(_02925_),
    .B(net3218),
    .Y(_02947_));
 sky130_fd_sc_hs__nor2_2 _08592_ (.A(net3171),
    .B(_02898_),
    .Y(_02948_));
 sky130_fd_sc_hs__nor3_1 _08593_ (.A(net3215),
    .B(net3221),
    .C(net3125),
    .Y(_02949_));
 sky130_fd_sc_hs__nand3_1 _08594_ (.A(net3606),
    .B(_00214_),
    .C(_00218_),
    .Y(_02950_));
 sky130_fd_sc_hs__and2_1 _08595_ (.A(_02911_),
    .B(_02900_),
    .X(_02951_));
 sky130_fd_sc_hs__inv_2 _08596_ (.A(_02951_),
    .Y(_02952_));
 sky130_fd_sc_hs__nor2_1 _08597_ (.A(net3216),
    .B(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hs__nor2_2 _08598_ (.A(net3296),
    .B(_02902_),
    .Y(_02954_));
 sky130_fd_sc_hs__nand3b_1 _08599_ (.A_N(net3261),
    .B(net3076),
    .C(net3257),
    .Y(_02955_));
 sky130_fd_sc_hs__nor2_1 _08600_ (.A(net3381),
    .B(_02955_),
    .Y(_02956_));
 sky130_fd_sc_hs__nand4_2 _08601_ (.A(net3077),
    .B(_02946_),
    .C(_02949_),
    .D(net2984),
    .Y(_02957_));
 sky130_fd_sc_hs__nor2_8 _08602_ (.A(_02957_),
    .B(net3131),
    .Y(_02958_));
 sky130_fd_sc_hs__nand2_2 _08603_ (.A(_02958_),
    .B(_02941_),
    .Y(_02959_));
 sky130_fd_sc_hs__nand2_1 _08604_ (.A(net3082),
    .B(_02881_),
    .Y(_02960_));
 sky130_fd_sc_hs__inv_1 _08605_ (.A(_02954_),
    .Y(_02961_));
 sky130_fd_sc_hs__nor3_1 _08606_ (.A(_02950_),
    .B(_02961_),
    .C(_02917_),
    .Y(_02962_));
 sky130_fd_sc_hs__nand2_1 _08607_ (.A(_02953_),
    .B(net3169),
    .Y(_02963_));
 sky130_fd_sc_hs__nor3_2 _08608_ (.A(_02947_),
    .B(_02898_),
    .C(_02963_),
    .Y(_02964_));
 sky130_fd_sc_hs__nor2_1 _08609_ (.A(_02929_),
    .B(net3221),
    .Y(_02965_));
 sky130_fd_sc_hs__nand3b_4 _08610_ (.A_N(net3125),
    .B(net2983),
    .C(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hs__nor3b_4 _08611_ (.A(_02960_),
    .B(_02966_),
    .C_N(net3078),
    .Y(_02967_));
 sky130_fd_sc_hs__nor2_1 _08612_ (.A(net3131),
    .B(_02967_),
    .Y(_02968_));
 sky130_fd_sc_hs__xor2_1 _08613_ (.A(_02968_),
    .B(net2987),
    .X(_02969_));
 sky130_fd_sc_hs__and2_2 _08614_ (.A(_02959_),
    .B(_02969_),
    .X(_02970_));
 sky130_fd_sc_hs__a21oi_1 _08615_ (.A1(net2987),
    .A2(net3084),
    .B1(net3131),
    .Y(_02971_));
 sky130_fd_sc_hs__nor2_1 _08616_ (.A(_02971_),
    .B(net2940),
    .Y(_02972_));
 sky130_fd_sc_hs__xnor2_1 _08617_ (.A(net3029),
    .B(_02972_),
    .Y(_02973_));
 sky130_fd_sc_hs__xor2_1 _08618_ (.A(net3084),
    .B(net2940),
    .X(_02974_));
 sky130_fd_sc_hs__nand3_2 _08619_ (.A(_02970_),
    .B(_02973_),
    .C(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hs__nand2_1 _08620_ (.A(net3606),
    .B(_00212_),
    .Y(_02976_));
 sky130_fd_sc_hs__nor3b_1 _08621_ (.A(_02976_),
    .B(net3213),
    .C_N(net3502),
    .Y(_02977_));
 sky130_fd_sc_hs__nand2_1 _08622_ (.A(net3176),
    .B(net3166),
    .Y(_02978_));
 sky130_fd_sc_hs__inv_1 _08623_ (.A(_02948_),
    .Y(_02979_));
 sky130_fd_sc_hs__nor3_4 _08624_ (.A(net3122),
    .B(net3124),
    .C(_02979_),
    .Y(_02980_));
 sky130_fd_sc_hs__nand4_2 _08625_ (.A(net2982),
    .B(net3168),
    .C(net3079),
    .D(net3081),
    .Y(_02981_));
 sky130_fd_sc_hs__o31ai_4 _08626_ (.A1(net2958),
    .A2(_02981_),
    .A3(net3028),
    .B1(net3086),
    .Y(_02982_));
 sky130_fd_sc_hs__xnor2_2 _08627_ (.A(_02982_),
    .B(net2989),
    .Y(_02983_));
 sky130_fd_sc_hs__nand2_1 _08628_ (.A(_02959_),
    .B(_02941_),
    .Y(_02984_));
 sky130_fd_sc_hs__nor2_1 _08629_ (.A(_02983_),
    .B(_02984_),
    .Y(_02985_));
 sky130_fd_sc_hs__nand2_2 _08630_ (.A(_02975_),
    .B(_02985_),
    .Y(_02986_));
 sky130_fd_sc_hs__nand2_2 _08631_ (.A(net2861),
    .B(net2888),
    .Y(_02987_));
 sky130_fd_sc_hs__nand2_2 _08632_ (.A(_02986_),
    .B(_02987_),
    .Y(_02988_));
 sky130_fd_sc_hs__nand3_2 _08633_ (.A(_02988_),
    .B(net2916),
    .C(net2851),
    .Y(_02989_));
 sky130_fd_sc_hs__a21oi_1 _08634_ (.A1(_02941_),
    .A2(net2888),
    .B1(net2887),
    .Y(_02990_));
 sky130_fd_sc_hs__nand2_1 _08635_ (.A(_02989_),
    .B(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hs__nand4_1 _08636_ (.A(net2939),
    .B(net3087),
    .C(net2990),
    .D(net2989),
    .Y(_02992_));
 sky130_fd_sc_hs__clkdlyinv3sd1_1 _08637_ (.A(net5127),
    .Y(_02993_));
 sky130_fd_sc_hs__a31oi_1 _08638_ (.A1(_02983_),
    .A2(_02969_),
    .A3(_02973_),
    .B1(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hs__or3_1 _08639_ (.A(net2958),
    .B(_02992_),
    .C(_02994_),
    .X(_02995_));
 sky130_fd_sc_hs__nand2_2 _08640_ (.A(_02991_),
    .B(_02995_),
    .Y(_02996_));
 sky130_fd_sc_hs__nand2_1 _08641_ (.A(_02988_),
    .B(net2916),
    .Y(_02997_));
 sky130_fd_sc_hs__inv_1 _08642_ (.A(net2916),
    .Y(_02998_));
 sky130_fd_sc_hs__nand3_1 _08643_ (.A(_02986_),
    .B(_02998_),
    .C(net2849),
    .Y(_02999_));
 sky130_fd_sc_hs__nand2_1 _08644_ (.A(net2956),
    .B(net3087),
    .Y(_03000_));
 sky130_fd_sc_hs__xnor2_1 _08645_ (.A(net3083),
    .B(_03000_),
    .Y(_03001_));
 sky130_fd_sc_hs__nand4_2 _08646_ (.A(_02997_),
    .B(_02999_),
    .C(_03001_),
    .D(net2851),
    .Y(_03002_));
 sky130_fd_sc_hs__or2b_1 _08647_ (.A(net2915),
    .B_N(_02986_),
    .X(_03003_));
 sky130_fd_sc_hs__nor2_1 _08648_ (.A(net2850),
    .B(_02988_),
    .Y(_03004_));
 sky130_fd_sc_hs__nor2_1 _08649_ (.A(_03003_),
    .B(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hs__nand3_2 _08650_ (.A(_03005_),
    .B(_03002_),
    .C(_02996_),
    .Y(_03006_));
 sky130_fd_sc_hs__inv_1 _08651_ (.A(net2802),
    .Y(_03007_));
 sky130_fd_sc_hs__nand2_2 _08652_ (.A(_03007_),
    .B(_03006_),
    .Y(_03008_));
 sky130_fd_sc_hs__nand2_2 _08653_ (.A(net2914),
    .B(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08654_ (.A(_03001_),
    .Y(_03010_));
 sky130_fd_sc_hs__nand3_2 _08655_ (.A(_03006_),
    .B(net2886),
    .C(_03007_),
    .Y(_03011_));
 sky130_fd_sc_hs__nand2_1 _08656_ (.A(net2959),
    .B(net3087),
    .Y(_03012_));
 sky130_fd_sc_hs__xnor2_1 _08657_ (.A(net3128),
    .B(_03012_),
    .Y(_03013_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08658_ (.A(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hs__nand2_1 _08659_ (.A(_02997_),
    .B(_02999_),
    .Y(_03015_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08660_ (.A(net2795),
    .Y(_03016_));
 sky130_fd_sc_hs__nand4_2 _08661_ (.A(_03009_),
    .B(_03011_),
    .C(_03014_),
    .D(_03016_),
    .Y(_03017_));
 sky130_fd_sc_hs__xnor2_2 _08662_ (.A(net2797),
    .B(net2791),
    .Y(_03018_));
 sky130_fd_sc_hs__nand2_1 _08663_ (.A(_03008_),
    .B(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08664_ (.A(net5168),
    .Y(_03020_));
 sky130_fd_sc_hs__nand3_1 _08665_ (.A(net2778),
    .B(net2796),
    .C(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hs__nand2_2 _08666_ (.A(_03019_),
    .B(_03021_),
    .Y(_03022_));
 sky130_fd_sc_hs__nor2_1 _08667_ (.A(_03010_),
    .B(_03015_),
    .Y(_03023_));
 sky130_fd_sc_hs__nand2b_1 _08668_ (.A_N(net2851),
    .B(_02997_),
    .Y(_03024_));
 sky130_fd_sc_hs__nand2_1 _08669_ (.A(_03024_),
    .B(net2803),
    .Y(_03025_));
 sky130_fd_sc_hs__xnor2_1 _08670_ (.A(_03023_),
    .B(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hs__nand2_1 _08671_ (.A(_03008_),
    .B(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hs__nand3b_1 _08672_ (.A_N(_03025_),
    .B(_03006_),
    .C(net2796),
    .Y(_03028_));
 sky130_fd_sc_hs__nand2_2 _08673_ (.A(_03027_),
    .B(_03028_),
    .Y(_03029_));
 sky130_fd_sc_hs__nor2_4 _08674_ (.A(_03022_),
    .B(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hs__nand2_2 _08675_ (.A(_03017_),
    .B(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hs__nand2_1 _08676_ (.A(net2792),
    .B(net2797),
    .Y(_03032_));
 sky130_fd_sc_hs__o21ai_1 _08677_ (.A1(_03007_),
    .A2(_03032_),
    .B1(net2806),
    .Y(_03033_));
 sky130_fd_sc_hs__nand2_1 _08678_ (.A(_03033_),
    .B(net2779),
    .Y(_03034_));
 sky130_fd_sc_hs__nand2_2 _08679_ (.A(_03031_),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hs__nand2_2 _08680_ (.A(net5129),
    .B(_03011_),
    .Y(_03036_));
 sky130_fd_sc_hs__nor2_4 _08681_ (.A(net2913),
    .B(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hs__a21oi_1 _08682_ (.A1(_03037_),
    .A2(net2790),
    .B1(net2754),
    .Y(_03038_));
 sky130_fd_sc_hs__nand2_2 _08683_ (.A(_03035_),
    .B(_03038_),
    .Y(_03039_));
 sky130_fd_sc_hs__nand2_1 _08684_ (.A(_03039_),
    .B(net2755),
    .Y(_03040_));
 sky130_fd_sc_hs__nand2_2 _08685_ (.A(_03040_),
    .B(net2738),
    .Y(_03041_));
 sky130_fd_sc_hs__nand2_2 _08686_ (.A(net2885),
    .B(_03035_),
    .Y(_03042_));
 sky130_fd_sc_hs__nand3_1 _08687_ (.A(_03031_),
    .B(net2913),
    .C(_03034_),
    .Y(_03043_));
 sky130_fd_sc_hs__nand2_1 _08688_ (.A(net2957),
    .B(net3088),
    .Y(_03044_));
 sky130_fd_sc_hs__xnor2_1 _08689_ (.A(net3126),
    .B(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hs__inv_1 _08690_ (.A(_03045_),
    .Y(_03046_));
 sky130_fd_sc_hs__and2_1 _08691_ (.A(net2761),
    .B(net2770),
    .X(_03047_));
 sky130_fd_sc_hs__nand4_2 _08692_ (.A(_03042_),
    .B(_03043_),
    .C(_03046_),
    .D(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hs__nand2_1 _08693_ (.A(net2760),
    .B(net2795),
    .Y(_03049_));
 sky130_fd_sc_hs__nand2_1 _08694_ (.A(net2771),
    .B(net2789),
    .Y(_03050_));
 sky130_fd_sc_hs__nand2_1 _08695_ (.A(_03049_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hs__xnor2_1 _08696_ (.A(_03051_),
    .B(_03037_),
    .Y(_03052_));
 sky130_fd_sc_hs__nand2_1 _08697_ (.A(_03035_),
    .B(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hs__nand3b_1 _08698_ (.A_N(_03051_),
    .B(_03031_),
    .C(_03034_),
    .Y(_03054_));
 sky130_fd_sc_hs__nand2_2 _08699_ (.A(_03053_),
    .B(_03054_),
    .Y(_03055_));
 sky130_fd_sc_hs__clkinv_1 _08700_ (.A(net2717),
    .Y(_03056_));
 sky130_fd_sc_hs__nand2_1 _08701_ (.A(net2718),
    .B(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hs__inv_1 _08702_ (.A(_03034_),
    .Y(_03058_));
 sky130_fd_sc_hs__o21ai_1 _08703_ (.A1(_03058_),
    .A2(net2748),
    .B1(net2756),
    .Y(_03059_));
 sky130_fd_sc_hs__nand2_1 _08704_ (.A(_03059_),
    .B(net2753),
    .Y(_03060_));
 sky130_fd_sc_hs__nand2_2 _08705_ (.A(_03039_),
    .B(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hs__o21ai_1 _08706_ (.A1(net2707),
    .A2(_03057_),
    .B1(net2716),
    .Y(_03062_));
 sky130_fd_sc_hs__nor2_2 _08707_ (.A(_03061_),
    .B(_03055_),
    .Y(_03063_));
 sky130_fd_sc_hs__nand2_2 _08708_ (.A(_03063_),
    .B(_03048_),
    .Y(_03064_));
 sky130_fd_sc_hs__nand2_2 _08709_ (.A(_03062_),
    .B(net2695),
    .Y(_03065_));
 sky130_fd_sc_hs__nand2_2 _08710_ (.A(_03041_),
    .B(_03064_),
    .Y(_03066_));
 sky130_fd_sc_hs__nand2_2 _08711_ (.A(net2884),
    .B(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hs__nand3_1 _08712_ (.A(_03064_),
    .B(net2912),
    .C(_03041_),
    .Y(_03068_));
 sky130_fd_sc_hs__a21oi_1 _08713_ (.A1(net3175),
    .A2(net3173),
    .B1(net3131),
    .Y(_03069_));
 sky130_fd_sc_hs__nor2_1 _08714_ (.A(net3131),
    .B(net2986),
    .Y(_03070_));
 sky130_fd_sc_hs__nor2_1 _08715_ (.A(_03069_),
    .B(_03070_),
    .Y(_03071_));
 sky130_fd_sc_hs__xnor2_1 _08716_ (.A(net3174),
    .B(_03071_),
    .Y(_03072_));
 sky130_fd_sc_hs__nand2_2 _08717_ (.A(_03042_),
    .B(_03043_),
    .Y(_03073_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08718_ (.A(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hs__nand4_2 _08719_ (.A(_03067_),
    .B(_03068_),
    .C(net2911),
    .D(_03074_),
    .Y(_03075_));
 sky130_fd_sc_hs__nand2_1 _08720_ (.A(_03042_),
    .B(net2752),
    .Y(_03076_));
 sky130_fd_sc_hs__nand2_1 _08721_ (.A(net2732),
    .B(net2747),
    .Y(_03077_));
 sky130_fd_sc_hs__nand2_1 _08722_ (.A(_03076_),
    .B(_03077_),
    .Y(_03078_));
 sky130_fd_sc_hs__nor2_2 _08723_ (.A(net2912),
    .B(_03073_),
    .Y(_03079_));
 sky130_fd_sc_hs__xnor2_1 _08724_ (.A(_03078_),
    .B(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hs__nand2_1 _08725_ (.A(_03080_),
    .B(_03066_),
    .Y(_03081_));
 sky130_fd_sc_hs__nand3b_1 _08726_ (.A_N(_03078_),
    .B(net5117),
    .C(_03041_),
    .Y(_03082_));
 sky130_fd_sc_hs__nand2_2 _08727_ (.A(_03081_),
    .B(_03082_),
    .Y(_03083_));
 sky130_fd_sc_hs__inv_1 _08728_ (.A(net2667),
    .Y(_03084_));
 sky130_fd_sc_hs__nand2_1 _08729_ (.A(net2669),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hs__nand3_1 _08730_ (.A(_03042_),
    .B(_03043_),
    .C(_03046_),
    .Y(_03086_));
 sky130_fd_sc_hs__nor2_1 _08731_ (.A(net2752),
    .B(_03086_),
    .Y(_03087_));
 sky130_fd_sc_hs__nand2_1 _08732_ (.A(_03087_),
    .B(net2717),
    .Y(_03088_));
 sky130_fd_sc_hs__nand2_1 _08733_ (.A(_03088_),
    .B(_03057_),
    .Y(_03089_));
 sky130_fd_sc_hs__nand2_1 _08734_ (.A(_03089_),
    .B(_03066_),
    .Y(_03090_));
 sky130_fd_sc_hs__nand3_1 _08735_ (.A(net5116),
    .B(_03041_),
    .C(net2717),
    .Y(_03091_));
 sky130_fd_sc_hs__nand2_2 _08736_ (.A(_03090_),
    .B(_03091_),
    .Y(_03092_));
 sky130_fd_sc_hs__o21ai_1 _08737_ (.A1(_03065_),
    .A2(_03085_),
    .B1(net2666),
    .Y(_03093_));
 sky130_fd_sc_hs__nor2_2 _08738_ (.A(_03083_),
    .B(_03092_),
    .Y(_03094_));
 sky130_fd_sc_hs__nand2_2 _08739_ (.A(_03094_),
    .B(_03075_),
    .Y(_03095_));
 sky130_fd_sc_hs__and2_2 _08740_ (.A(_03093_),
    .B(net2648),
    .X(_03096_));
 sky130_fd_sc_hs__nand2_2 _08741_ (.A(_03095_),
    .B(_03065_),
    .Y(_03097_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08742_ (.A(_03072_),
    .Y(_03098_));
 sky130_fd_sc_hs__nand2_2 _08743_ (.A(_03067_),
    .B(_03068_),
    .Y(_03099_));
 sky130_fd_sc_hs__nor3_2 _08744_ (.A(_03098_),
    .B(net2715),
    .C(_03099_),
    .Y(_03100_));
 sky130_fd_sc_hs__nor2_1 _08745_ (.A(net2668),
    .B(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hs__nand2_2 _08746_ (.A(_03097_),
    .B(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hs__o21ai_1 _08747_ (.A1(_03065_),
    .A2(_03100_),
    .B1(net2668),
    .Y(_03103_));
 sky130_fd_sc_hs__nand2_2 _08748_ (.A(_03102_),
    .B(_03103_),
    .Y(_03104_));
 sky130_fd_sc_hs__nand2_1 _08749_ (.A(net2673),
    .B(net2715),
    .Y(_03105_));
 sky130_fd_sc_hs__nand2_1 _08750_ (.A(net2688),
    .B(net2706),
    .Y(_03106_));
 sky130_fd_sc_hs__nand2_1 _08751_ (.A(_03105_),
    .B(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hs__nor2_2 _08752_ (.A(_03098_),
    .B(_03099_),
    .Y(_03108_));
 sky130_fd_sc_hs__xnor2_2 _08753_ (.A(_03107_),
    .B(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hs__nand2_2 _08754_ (.A(_03109_),
    .B(_03097_),
    .Y(_03110_));
 sky130_fd_sc_hs__nand3b_1 _08755_ (.A_N(_03107_),
    .B(net2648),
    .C(net2675),
    .Y(_03111_));
 sky130_fd_sc_hs__nand2_2 _08756_ (.A(_03111_),
    .B(_03110_),
    .Y(_03112_));
 sky130_fd_sc_hs__nor2_4 _08757_ (.A(_03104_),
    .B(_03112_),
    .Y(_03113_));
 sky130_fd_sc_hs__nand2_2 _08758_ (.A(net2911),
    .B(_03097_),
    .Y(_03114_));
 sky130_fd_sc_hs__nand3_1 _08759_ (.A(_03095_),
    .B(net2883),
    .C(net2674),
    .Y(_03115_));
 sky130_fd_sc_hs__nand2_1 _08760_ (.A(net2982),
    .B(net3168),
    .Y(_03116_));
 sky130_fd_sc_hs__nand2_1 _08761_ (.A(_03116_),
    .B(net3088),
    .Y(_03117_));
 sky130_fd_sc_hs__xnor2_1 _08762_ (.A(net3173),
    .B(_03117_),
    .Y(_03118_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08763_ (.A(net2665),
    .Y(_03119_));
 sky130_fd_sc_hs__nand4_2 _08764_ (.A(_03114_),
    .B(_03115_),
    .C(net2910),
    .D(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hs__o21ai_1 _08765_ (.A1(net2631),
    .A2(_03113_),
    .B1(net5110),
    .Y(_03121_));
 sky130_fd_sc_hs__nand2_1 _08766_ (.A(net2624),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hs__and2_1 _08767_ (.A(_03102_),
    .B(_03103_),
    .X(_03123_));
 sky130_fd_sc_hs__inv_1 _08768_ (.A(_03112_),
    .Y(_03124_));
 sky130_fd_sc_hs__o211ai_1 _08769_ (.A1(_03123_),
    .A2(_03096_),
    .B1(_03124_),
    .C1(net5112),
    .Y(_03125_));
 sky130_fd_sc_hs__and2_1 _08770_ (.A(_03122_),
    .B(_03125_),
    .X(_03126_));
 sky130_fd_sc_hs__bufinv_8 _08771_ (.A(_03096_),
    .Y(_03127_));
 sky130_fd_sc_hs__nand2_1 _08772_ (.A(net5111),
    .B(_03124_),
    .Y(_03128_));
 sky130_fd_sc_hs__o21ai_1 _08773_ (.A1(_03127_),
    .A2(_03128_),
    .B1(net2625),
    .Y(_03129_));
 sky130_fd_sc_hs__nand2_2 _08774_ (.A(_03120_),
    .B(_03113_),
    .Y(_03130_));
 sky130_fd_sc_hs__and2_2 _08775_ (.A(net2612),
    .B(_03129_),
    .X(_03131_));
 sky130_fd_sc_hs__nand2_1 _08776_ (.A(_03114_),
    .B(net2665),
    .Y(_03132_));
 sky130_fd_sc_hs__nand2_1 _08777_ (.A(net2642),
    .B(net2660),
    .Y(_03133_));
 sky130_fd_sc_hs__nand2_1 _08778_ (.A(_03132_),
    .B(_03133_),
    .Y(_03134_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08779_ (.A(net2910),
    .Y(_03135_));
 sky130_fd_sc_hs__nand2_1 _08780_ (.A(net2630),
    .B(net2641),
    .Y(_03136_));
 sky130_fd_sc_hs__nor2_2 _08781_ (.A(_03135_),
    .B(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hs__xnor2_1 _08782_ (.A(_03134_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hs__nand2_2 _08783_ (.A(_03130_),
    .B(_03127_),
    .Y(_03139_));
 sky130_fd_sc_hs__nand2_1 _08784_ (.A(_03138_),
    .B(_03139_),
    .Y(_03140_));
 sky130_fd_sc_hs__inv_1 _08785_ (.A(_03134_),
    .Y(_03141_));
 sky130_fd_sc_hs__nand3_1 _08786_ (.A(_03130_),
    .B(_03127_),
    .C(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hs__nand2_2 _08787_ (.A(_03140_),
    .B(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hs__inv_1 _08788_ (.A(_03143_),
    .Y(_03144_));
 sky130_fd_sc_hs__nand3_2 _08789_ (.A(_03130_),
    .B(net2910),
    .C(_03127_),
    .Y(_03145_));
 sky130_fd_sc_hs__o21ai_1 _08790_ (.A1(net2631),
    .A2(_03113_),
    .B1(net2882),
    .Y(_03146_));
 sky130_fd_sc_hs__nand2_2 _08791_ (.A(_03146_),
    .B(_03145_),
    .Y(_03147_));
 sky130_fd_sc_hs__xnor2_1 _08792_ (.A(net3214),
    .B(net2955),
    .Y(_03148_));
 sky130_fd_sc_hs__inv_1 _08793_ (.A(net2623),
    .Y(_03149_));
 sky130_fd_sc_hs__nand3_4 _08794_ (.A(_03147_),
    .B(net2938),
    .C(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hs__o211ai_1 _08795_ (.A1(_03126_),
    .A2(_03131_),
    .B1(net2576),
    .C1(net2587),
    .Y(_03151_));
 sky130_fd_sc_hs__a21o_1 _08796_ (.A1(net2587),
    .A2(_03131_),
    .B1(_03144_),
    .X(_03152_));
 sky130_fd_sc_hs__and2_1 _08797_ (.A(_03151_),
    .B(_03152_),
    .X(_03153_));
 sky130_fd_sc_hs__inv_4 _08798_ (.A(_03131_),
    .Y(_03154_));
 sky130_fd_sc_hs__nand2_1 _08799_ (.A(_03144_),
    .B(_03150_),
    .Y(_03155_));
 sky130_fd_sc_hs__nand2_2 _08800_ (.A(_03122_),
    .B(_03125_),
    .Y(_03156_));
 sky130_fd_sc_hs__o21ai_2 _08801_ (.A1(_03154_),
    .A2(_03155_),
    .B1(net2592),
    .Y(_03157_));
 sky130_fd_sc_hs__nor2_4 _08802_ (.A(_03143_),
    .B(_03156_),
    .Y(_03158_));
 sky130_fd_sc_hs__nand2_2 _08803_ (.A(_03150_),
    .B(_03158_),
    .Y(_03159_));
 sky130_fd_sc_hs__and2_2 _08804_ (.A(_03159_),
    .B(_03157_),
    .X(_03160_));
 sky130_fd_sc_hs__nand2_2 _08805_ (.A(_03154_),
    .B(_03159_),
    .Y(_03161_));
 sky130_fd_sc_hs__xnor2_1 _08806_ (.A(net2910),
    .B(net2623),
    .Y(_03162_));
 sky130_fd_sc_hs__nand2_1 _08807_ (.A(net2603),
    .B(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hs__o21ai_2 _08808_ (.A1(net2623),
    .A2(net2603),
    .B1(_03163_),
    .Y(_03164_));
 sky130_fd_sc_hs__nand2_1 _08809_ (.A(_03147_),
    .B(net2938),
    .Y(_03165_));
 sky130_fd_sc_hs__xnor2_1 _08810_ (.A(_03164_),
    .B(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hs__nand2_1 _08811_ (.A(_03161_),
    .B(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hs__nand3_1 _08812_ (.A(_03159_),
    .B(_03154_),
    .C(_03164_),
    .Y(_03168_));
 sky130_fd_sc_hs__nand2_2 _08813_ (.A(_03167_),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hs__inv_1 _08814_ (.A(net5179),
    .Y(_03170_));
 sky130_fd_sc_hs__nand2_2 _08815_ (.A(_03161_),
    .B(net2938),
    .Y(_03171_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08816_ (.A(net2938),
    .Y(_03172_));
 sky130_fd_sc_hs__nand3_2 _08817_ (.A(net5173),
    .B(_03172_),
    .C(_03154_),
    .Y(_03173_));
 sky130_fd_sc_hs__or2_1 _08818_ (.A(net3132),
    .B(net2983),
    .X(_03174_));
 sky130_fd_sc_hs__xnor2_1 _08819_ (.A(net3221),
    .B(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08820_ (.A(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hs__nand4_2 _08821_ (.A(_03173_),
    .B(_03171_),
    .C(_03176_),
    .D(net2593),
    .Y(_03177_));
 sky130_fd_sc_hs__o211ai_1 _08822_ (.A1(_03153_),
    .A2(net2550),
    .B1(_03170_),
    .C1(net5122),
    .Y(_03178_));
 sky130_fd_sc_hs__nand2_2 _08823_ (.A(_03151_),
    .B(_03152_),
    .Y(_03179_));
 sky130_fd_sc_hs__nand2_1 _08824_ (.A(_03178_),
    .B(net2560),
    .Y(_03180_));
 sky130_fd_sc_hs__nor2_4 _08825_ (.A(_03169_),
    .B(_03179_),
    .Y(_03181_));
 sky130_fd_sc_hs__nand2_2 _08826_ (.A(_03181_),
    .B(_03177_),
    .Y(_03182_));
 sky130_fd_sc_hs__and2_1 _08827_ (.A(_03180_),
    .B(net5114),
    .X(_03183_));
 sky130_fd_sc_hs__bufinv_8 _08828_ (.A(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hs__nand2_1 _08829_ (.A(net2548),
    .B(net2561),
    .Y(_03185_));
 sky130_fd_sc_hs__bufinv_8 _08830_ (.A(_03160_),
    .Y(_03186_));
 sky130_fd_sc_hs__nand3_2 _08831_ (.A(_03182_),
    .B(_03176_),
    .C(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hs__o21ai_1 _08832_ (.A1(net2549),
    .A2(net5134),
    .B1(_03175_),
    .Y(_03188_));
 sky130_fd_sc_hs__nand2_2 _08833_ (.A(_03188_),
    .B(_03187_),
    .Y(_03189_));
 sky130_fd_sc_hs__a31o_1 _08834_ (.A1(net3080),
    .A2(net3220),
    .A3(net3259),
    .B1(net3132),
    .X(_03190_));
 sky130_fd_sc_hs__xnor2_1 _08835_ (.A(net3177),
    .B(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hs__nand2_1 _08836_ (.A(net2507),
    .B(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hs__nand2_2 _08837_ (.A(_03182_),
    .B(_03186_),
    .Y(_03193_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08838_ (.A(net2593),
    .Y(_03194_));
 sky130_fd_sc_hs__nand2_1 _08839_ (.A(_03171_),
    .B(_03194_),
    .Y(_03195_));
 sky130_fd_sc_hs__nand3_1 _08840_ (.A(net5180),
    .B(net2938),
    .C(net2593),
    .Y(_03196_));
 sky130_fd_sc_hs__and2_2 _08841_ (.A(_03195_),
    .B(_03196_),
    .X(_03197_));
 sky130_fd_sc_hs__nand3_1 _08842_ (.A(net2548),
    .B(net2561),
    .C(_03176_),
    .Y(_03198_));
 sky130_fd_sc_hs__nand2_1 _08843_ (.A(_03197_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hs__nand4_1 _08844_ (.A(net2548),
    .B(net2561),
    .C(_03176_),
    .D(net2586),
    .Y(_03200_));
 sky130_fd_sc_hs__nand2_1 _08845_ (.A(_03199_),
    .B(_03200_),
    .Y(_03201_));
 sky130_fd_sc_hs__nand2_1 _08846_ (.A(_03193_),
    .B(_03201_),
    .Y(_03202_));
 sky130_fd_sc_hs__nand3_1 _08847_ (.A(_03182_),
    .B(_03197_),
    .C(_03186_),
    .Y(_03203_));
 sky130_fd_sc_hs__nand2_2 _08848_ (.A(_03203_),
    .B(_03202_),
    .Y(_03204_));
 sky130_fd_sc_hs__o21bai_1 _08849_ (.A1(net2542),
    .A2(_03192_),
    .B1_N(net5182),
    .Y(_03205_));
 sky130_fd_sc_hs__o21ai_1 _08850_ (.A1(_03160_),
    .A2(_03181_),
    .B1(net5122),
    .Y(_03206_));
 sky130_fd_sc_hs__nand2_1 _08851_ (.A(_03206_),
    .B(net2543),
    .Y(_03207_));
 sky130_fd_sc_hs__nand2_1 _08852_ (.A(_03178_),
    .B(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hs__o21ai_2 _08853_ (.A1(_03184_),
    .A2(_03205_),
    .B1(net2506),
    .Y(_03209_));
 sky130_fd_sc_hs__clkinv_1 _08854_ (.A(_03185_),
    .Y(_03210_));
 sky130_fd_sc_hs__nand3_2 _08855_ (.A(_03210_),
    .B(_03191_),
    .C(_03189_),
    .Y(_03211_));
 sky130_fd_sc_hs__nor2_4 _08856_ (.A(_03204_),
    .B(_03208_),
    .Y(_03212_));
 sky130_fd_sc_hs__nand2_2 _08857_ (.A(_03211_),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hs__and2_1 _08858_ (.A(_03209_),
    .B(net2485),
    .X(_03214_));
 sky130_fd_sc_hs__nand2_8 _08859_ (.A(_03213_),
    .B(_03184_),
    .Y(_03215_));
 sky130_fd_sc_hs__xnor2_1 _08860_ (.A(_03176_),
    .B(_03185_),
    .Y(_03216_));
 sky130_fd_sc_hs__nand2_1 _08861_ (.A(net2518),
    .B(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hs__nand3_1 _08862_ (.A(net2526),
    .B(_03210_),
    .C(net2541),
    .Y(_03218_));
 sky130_fd_sc_hs__nand4_1 _08863_ (.A(_03189_),
    .B(_03191_),
    .C(_03217_),
    .D(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hs__o21ai_1 _08864_ (.A1(net2542),
    .A2(net2518),
    .B1(_03217_),
    .Y(_03220_));
 sky130_fd_sc_hs__nand2_1 _08865_ (.A(_03192_),
    .B(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hs__nand2_1 _08866_ (.A(_03219_),
    .B(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hs__nand2_2 _08867_ (.A(_03215_),
    .B(_03222_),
    .Y(_03223_));
 sky130_fd_sc_hs__nand3_1 _08868_ (.A(_03213_),
    .B(_03220_),
    .C(_03184_),
    .Y(_03224_));
 sky130_fd_sc_hs__nand2_2 _08869_ (.A(_03223_),
    .B(_03224_),
    .Y(_03225_));
 sky130_fd_sc_hs__o21ai_1 _08870_ (.A1(net2509),
    .A2(net2490),
    .B1(net2497),
    .Y(_03226_));
 sky130_fd_sc_hs__nand2_1 _08871_ (.A(_03226_),
    .B(net2499),
    .Y(_03227_));
 sky130_fd_sc_hs__a31oi_2 _08872_ (.A1(net2507),
    .A2(_03191_),
    .A3(net2532),
    .B1(net2498),
    .Y(_03228_));
 sky130_fd_sc_hs__nand2_2 _08873_ (.A(_03228_),
    .B(_03215_),
    .Y(_03229_));
 sky130_fd_sc_hs__nand2_2 _08874_ (.A(_03229_),
    .B(_03227_),
    .Y(_03230_));
 sky130_fd_sc_hs__nor2_4 _08875_ (.A(_03230_),
    .B(_03225_),
    .Y(_03231_));
 sky130_fd_sc_hs__nand2_2 _08876_ (.A(_03215_),
    .B(_03191_),
    .Y(_03232_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08877_ (.A(_03191_),
    .Y(_03233_));
 sky130_fd_sc_hs__nand3_2 _08878_ (.A(net5167),
    .B(_03233_),
    .C(_03184_),
    .Y(_03234_));
 sky130_fd_sc_hs__o31ai_1 _08879_ (.A1(net3123),
    .A2(net3172),
    .A3(net3124),
    .B1(net3089),
    .Y(_03235_));
 sky130_fd_sc_hs__xnor2_1 _08880_ (.A(net3220),
    .B(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hs__nand4_2 _08881_ (.A(_03232_),
    .B(_03234_),
    .C(_03236_),
    .D(net2508),
    .Y(_03237_));
 sky130_fd_sc_hs__o21ai_2 _08882_ (.A1(_03214_),
    .A2(net2446),
    .B1(net2456),
    .Y(_03238_));
 sky130_fd_sc_hs__nand2_2 _08883_ (.A(_03238_),
    .B(net2458),
    .Y(_03239_));
 sky130_fd_sc_hs__nand2_2 _08884_ (.A(_03237_),
    .B(_03231_),
    .Y(_03240_));
 sky130_fd_sc_hs__nand2_1 _08885_ (.A(_03209_),
    .B(net2485),
    .Y(_03241_));
 sky130_fd_sc_hs__nand2_8 _08886_ (.A(net2474),
    .B(_03240_),
    .Y(_03242_));
 sky130_fd_sc_hs__and2_1 _08887_ (.A(_03223_),
    .B(net2477),
    .X(_03243_));
 sky130_fd_sc_hs__and2_1 _08888_ (.A(_03237_),
    .B(_03243_),
    .X(_03244_));
 sky130_fd_sc_hs__nand2_2 _08889_ (.A(_03244_),
    .B(_03242_),
    .Y(_03245_));
 sky130_fd_sc_hs__and2_2 _08890_ (.A(_03239_),
    .B(net5138),
    .X(_03246_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08891_ (.A(net2508),
    .Y(_03247_));
 sky130_fd_sc_hs__xnor2_1 _08892_ (.A(_03233_),
    .B(net2508),
    .Y(_03248_));
 sky130_fd_sc_hs__nand2_1 _08893_ (.A(net5137),
    .B(_03248_),
    .Y(_03249_));
 sky130_fd_sc_hs__o21ai_4 _08894_ (.A1(_03247_),
    .A2(net5137),
    .B1(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hs__nand3_2 _08895_ (.A(net2463),
    .B(net2476),
    .C(_03236_),
    .Y(_03251_));
 sky130_fd_sc_hs__xor2_1 _08896_ (.A(_03250_),
    .B(net2454),
    .X(_03252_));
 sky130_fd_sc_hs__nand2_1 _08897_ (.A(_03252_),
    .B(_03242_),
    .Y(_03253_));
 sky130_fd_sc_hs__nand3b_1 _08898_ (.A_N(net2455),
    .B(net2436),
    .C(net2475),
    .Y(_03254_));
 sky130_fd_sc_hs__nand2_2 _08899_ (.A(_03253_),
    .B(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hs__nand2_8 _08900_ (.A(_03242_),
    .B(_03236_),
    .Y(_03256_));
 sky130_fd_sc_hs__and2_1 _08901_ (.A(net5171),
    .B(net5178),
    .X(_03257_));
 sky130_fd_sc_hs__nand2_1 _08902_ (.A(_03257_),
    .B(_03243_),
    .Y(_03258_));
 sky130_fd_sc_hs__inv_1 _08903_ (.A(_03236_),
    .Y(_03259_));
 sky130_fd_sc_hs__nand3_1 _08904_ (.A(_03258_),
    .B(_03259_),
    .C(net2474),
    .Y(_03260_));
 sky130_fd_sc_hs__and2_1 _08905_ (.A(net2463),
    .B(net2476),
    .X(_03261_));
 sky130_fd_sc_hs__and2_1 _08906_ (.A(_03260_),
    .B(_03261_),
    .X(_03262_));
 sky130_fd_sc_hs__nand2_8 _08907_ (.A(_03262_),
    .B(_03256_),
    .Y(_03263_));
 sky130_fd_sc_hs__nand3_2 _08908_ (.A(_03246_),
    .B(_03255_),
    .C(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hs__nand2_1 _08909_ (.A(_03245_),
    .B(net2457),
    .Y(_03265_));
 sky130_fd_sc_hs__nand2_1 _08910_ (.A(_03265_),
    .B(net2437),
    .Y(_03266_));
 sky130_fd_sc_hs__nand2_2 _08911_ (.A(_03264_),
    .B(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hs__or2_1 _08912_ (.A(net3080),
    .B(net3132),
    .X(_03268_));
 sky130_fd_sc_hs__xnor2_1 _08913_ (.A(net3259),
    .B(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hs__nand2_2 _08914_ (.A(_03267_),
    .B(_03269_),
    .Y(_03270_));
 sky130_fd_sc_hs__xnor2_1 _08915_ (.A(_03250_),
    .B(_03251_),
    .Y(_03271_));
 sky130_fd_sc_hs__nand2_2 _08916_ (.A(_03242_),
    .B(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hs__nand3_4 _08917_ (.A(net2436),
    .B(net2475),
    .C(net2455),
    .Y(_03273_));
 sky130_fd_sc_hs__nand2_8 _08918_ (.A(_03273_),
    .B(_03272_),
    .Y(_03274_));
 sky130_fd_sc_hs__nand2_2 _08919_ (.A(_03245_),
    .B(_03239_),
    .Y(_03275_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08920_ (.A(_03269_),
    .Y(_03276_));
 sky130_fd_sc_hs__o211ai_2 _08921_ (.A1(net5181),
    .A2(net5142),
    .B1(_03276_),
    .C1(_03266_),
    .Y(_03277_));
 sky130_fd_sc_hs__nand2_1 _08922_ (.A(net3027),
    .B(net3089),
    .Y(_03278_));
 sky130_fd_sc_hs__xnor2_1 _08923_ (.A(net3219),
    .B(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hs__and2_2 _08924_ (.A(_03256_),
    .B(net2435),
    .X(_03280_));
 sky130_fd_sc_hs__nand4_2 _08925_ (.A(_03277_),
    .B(_03270_),
    .C(net2954),
    .D(net2401),
    .Y(_03281_));
 sky130_fd_sc_hs__nor2_8 _08926_ (.A(_03275_),
    .B(_03274_),
    .Y(_03282_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08927_ (.A(net2954),
    .Y(_03283_));
 sky130_fd_sc_hs__nand2_1 _08928_ (.A(_03283_),
    .B(_03276_),
    .Y(_03284_));
 sky130_fd_sc_hs__nand3_1 _08929_ (.A(net2415),
    .B(net2429),
    .C(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hs__nand2_1 _08930_ (.A(_03282_),
    .B(_03285_),
    .Y(_03286_));
 sky130_fd_sc_hs__nand2_1 _08931_ (.A(_03276_),
    .B(net2954),
    .Y(_03287_));
 sky130_fd_sc_hs__nor2_2 _08932_ (.A(_03287_),
    .B(_03263_),
    .Y(_03288_));
 sky130_fd_sc_hs__nand2_2 _08933_ (.A(_03282_),
    .B(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hs__nand3_2 _08934_ (.A(_03289_),
    .B(_03286_),
    .C(_03266_),
    .Y(_03290_));
 sky130_fd_sc_hs__xnor2_2 _08935_ (.A(net2453),
    .B(_03256_),
    .Y(_03291_));
 sky130_fd_sc_hs__nand2_1 _08936_ (.A(_03280_),
    .B(_03269_),
    .Y(_03292_));
 sky130_fd_sc_hs__nand2_1 _08937_ (.A(_03291_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hs__inv_1 _08938_ (.A(net2453),
    .Y(_03294_));
 sky130_fd_sc_hs__nand4_1 _08939_ (.A(net2416),
    .B(_03269_),
    .C(_03294_),
    .D(net2435),
    .Y(_03295_));
 sky130_fd_sc_hs__nand2_2 _08940_ (.A(_03293_),
    .B(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hs__nand2_2 _08941_ (.A(_03296_),
    .B(_03290_),
    .Y(_03297_));
 sky130_fd_sc_hs__and2_2 _08942_ (.A(_03264_),
    .B(_03266_),
    .X(_03298_));
 sky130_fd_sc_hs__inv_1 _08943_ (.A(_03263_),
    .Y(_03299_));
 sky130_fd_sc_hs__nand3_1 _08944_ (.A(_03282_),
    .B(_03299_),
    .C(_03276_),
    .Y(_03300_));
 sky130_fd_sc_hs__nand3_2 _08945_ (.A(_03298_),
    .B(_03291_),
    .C(_03300_),
    .Y(_03301_));
 sky130_fd_sc_hs__and2_2 _08946_ (.A(_03297_),
    .B(_03301_),
    .X(_03302_));
 sky130_fd_sc_hs__a21boi_1 _08947_ (.A1(net5138),
    .A2(net2457),
    .B1_N(net2437),
    .Y(_03303_));
 sky130_fd_sc_hs__o22ai_1 _08948_ (.A1(_03276_),
    .A2(net5108),
    .B1(_03303_),
    .B2(net2394),
    .Y(_03304_));
 sky130_fd_sc_hs__nand2_1 _08949_ (.A(_03304_),
    .B(net2404),
    .Y(_03305_));
 sky130_fd_sc_hs__o211ai_1 _08950_ (.A1(_03276_),
    .A2(_03263_),
    .B1(_03274_),
    .C1(_03303_),
    .Y(_03306_));
 sky130_fd_sc_hs__nand2_1 _08951_ (.A(_03305_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hs__nand3_2 _08952_ (.A(_03281_),
    .B(_03302_),
    .C(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hs__nor2_2 _08953_ (.A(_03276_),
    .B(_03263_),
    .Y(_03309_));
 sky130_fd_sc_hs__nor2_2 _08954_ (.A(net2403),
    .B(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hs__nand2_2 _08955_ (.A(_03290_),
    .B(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hs__nand2_1 _08956_ (.A(_03311_),
    .B(net2402),
    .Y(_03312_));
 sky130_fd_sc_hs__nand2_1 _08957_ (.A(_03310_),
    .B(net2405),
    .Y(_03313_));
 sky130_fd_sc_hs__nand2_1 _08958_ (.A(_03312_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hs__nand2_2 _08959_ (.A(_03314_),
    .B(_03308_),
    .Y(_03315_));
 sky130_fd_sc_hs__and2_1 _08960_ (.A(net2380),
    .B(net2388),
    .X(_03316_));
 sky130_fd_sc_hs__nand3_1 _08961_ (.A(_03315_),
    .B(net2954),
    .C(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hs__xor2_1 _08962_ (.A(net2401),
    .B(net2380),
    .X(_03318_));
 sky130_fd_sc_hs__nand2_1 _08963_ (.A(_03317_),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hs__inv_2 _08964_ (.A(net2365),
    .Y(_03320_));
 sky130_fd_sc_hs__nand2_1 _08965_ (.A(_03315_),
    .B(net2356),
    .Y(_03321_));
 sky130_fd_sc_hs__nand2_1 _08966_ (.A(_03319_),
    .B(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hs__nand3_2 _08967_ (.A(_03314_),
    .B(net2954),
    .C(_03308_),
    .Y(_03323_));
 sky130_fd_sc_hs__and2_2 _08968_ (.A(_03312_),
    .B(_03313_),
    .X(_03324_));
 sky130_fd_sc_hs__xnor2_1 _08969_ (.A(net2403),
    .B(net2393),
    .Y(_03325_));
 sky130_fd_sc_hs__nand2_1 _08970_ (.A(net2379),
    .B(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hs__nand3_1 _08971_ (.A(net2387),
    .B(net2403),
    .C(net2386),
    .Y(_03327_));
 sky130_fd_sc_hs__nand2_2 _08972_ (.A(_03327_),
    .B(_03326_),
    .Y(_03328_));
 sky130_fd_sc_hs__nand2_2 _08973_ (.A(net2364),
    .B(net2378),
    .Y(_03329_));
 sky130_fd_sc_hs__nor2_4 _08974_ (.A(_03328_),
    .B(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hs__o21ai_4 _08975_ (.A1(_03330_),
    .A2(_03324_),
    .B1(_03283_),
    .Y(_03331_));
 sky130_fd_sc_hs__nand2_2 _08976_ (.A(_03331_),
    .B(_03323_),
    .Y(_03332_));
 sky130_fd_sc_hs__nand2_1 _08977_ (.A(net3089),
    .B(net3127),
    .Y(_03333_));
 sky130_fd_sc_hs__xnor2_1 _08978_ (.A(net3297),
    .B(_03333_),
    .Y(_03334_));
 sky130_fd_sc_hs__nand3_2 _08979_ (.A(net2363),
    .B(_03334_),
    .C(_03332_),
    .Y(_03335_));
 sky130_fd_sc_hs__xnor2_1 _08980_ (.A(net2365),
    .B(net2357),
    .Y(_03336_));
 sky130_fd_sc_hs__nand2_1 _08981_ (.A(_03315_),
    .B(_03336_),
    .Y(_03337_));
 sky130_fd_sc_hs__o21a_2 _08982_ (.A1(net2357),
    .A2(_03315_),
    .B1(_03337_),
    .X(_03338_));
 sky130_fd_sc_hs__nand3_2 _08983_ (.A(_03338_),
    .B(_03322_),
    .C(_03335_),
    .Y(_03339_));
 sky130_fd_sc_hs__o31ai_1 _08984_ (.A1(_03329_),
    .A2(_03320_),
    .A3(_03314_),
    .B1(net2355),
    .Y(_03340_));
 sky130_fd_sc_hs__nand2_1 _08985_ (.A(_03340_),
    .B(net2351),
    .Y(_03341_));
 sky130_fd_sc_hs__nand2_2 _08986_ (.A(net2329),
    .B(_03339_),
    .Y(_03342_));
 sky130_fd_sc_hs__nand2_2 _08987_ (.A(_03342_),
    .B(_03334_),
    .Y(_03343_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _08988_ (.A(_03334_),
    .Y(_03344_));
 sky130_fd_sc_hs__nand3_2 _08989_ (.A(net5177),
    .B(_03344_),
    .C(net2329),
    .Y(_03345_));
 sky130_fd_sc_hs__nand2_1 _08990_ (.A(net3089),
    .B(net3123),
    .Y(_03346_));
 sky130_fd_sc_hs__xnor2_1 _08991_ (.A(net3217),
    .B(_03346_),
    .Y(_03347_));
 sky130_fd_sc_hs__nand4_2 _08992_ (.A(_03345_),
    .B(_03343_),
    .C(_03347_),
    .D(net2331),
    .Y(_03348_));
 sky130_fd_sc_hs__and2_2 _08993_ (.A(net2321),
    .B(net2332),
    .X(_03349_));
 sky130_fd_sc_hs__nand2_1 _08994_ (.A(net2330),
    .B(net2363),
    .Y(_03350_));
 sky130_fd_sc_hs__nor2_1 _08995_ (.A(_03344_),
    .B(_03350_),
    .Y(_03351_));
 sky130_fd_sc_hs__nand2_1 _08996_ (.A(_03349_),
    .B(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hs__nand2_1 _08997_ (.A(net2311),
    .B(net2320),
    .Y(_03353_));
 sky130_fd_sc_hs__nand2_2 _08998_ (.A(_03352_),
    .B(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hs__nand2_1 _08999_ (.A(_03342_),
    .B(_03354_),
    .Y(_03355_));
 sky130_fd_sc_hs__nand3_1 _09000_ (.A(net2305),
    .B(_03349_),
    .C(net2329),
    .Y(_03356_));
 sky130_fd_sc_hs__nand2_2 _09001_ (.A(_03355_),
    .B(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hs__a21oi_1 _09002_ (.A1(net2342),
    .A2(net2341),
    .B1(_03344_),
    .Y(_03358_));
 sky130_fd_sc_hs__nand2_1 _09003_ (.A(net2343),
    .B(net2954),
    .Y(_03359_));
 sky130_fd_sc_hs__xor2_2 _09004_ (.A(_03359_),
    .B(net2363),
    .X(_03360_));
 sky130_fd_sc_hs__xnor2_1 _09005_ (.A(_03358_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hs__nand2_2 _09006_ (.A(_03361_),
    .B(_03342_),
    .Y(_03362_));
 sky130_fd_sc_hs__nand3b_1 _09007_ (.A_N(_03360_),
    .B(_03339_),
    .C(net2329),
    .Y(_03363_));
 sky130_fd_sc_hs__nand2_2 _09008_ (.A(_03363_),
    .B(_03362_),
    .Y(_03364_));
 sky130_fd_sc_hs__nor2_4 _09009_ (.A(_03364_),
    .B(_03357_),
    .Y(_03365_));
 sky130_fd_sc_hs__nand2_2 _09010_ (.A(_03365_),
    .B(_03348_),
    .Y(_03366_));
 sky130_fd_sc_hs__or3_1 _09011_ (.A(net2319),
    .B(net2329),
    .C(_03353_),
    .X(_03367_));
 sky130_fd_sc_hs__o21ai_1 _09012_ (.A1(net2310),
    .A2(_03349_),
    .B1(net2319),
    .Y(_03368_));
 sky130_fd_sc_hs__nand2_2 _09013_ (.A(_03367_),
    .B(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hs__inv_2 _09014_ (.A(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hs__nand2_2 _09015_ (.A(_03370_),
    .B(_03366_),
    .Y(_03371_));
 sky130_fd_sc_hs__nand2_2 _09016_ (.A(_03371_),
    .B(_03347_),
    .Y(_03372_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09017_ (.A(_03347_),
    .Y(_03373_));
 sky130_fd_sc_hs__nand3_2 _09018_ (.A(net5140),
    .B(_03373_),
    .C(_03370_),
    .Y(_03374_));
 sky130_fd_sc_hs__o31ai_1 _09019_ (.A1(_02909_),
    .A2(net3261),
    .A3(net3293),
    .B1(net3089),
    .Y(_03375_));
 sky130_fd_sc_hs__xnor2_1 _09020_ (.A(net3332),
    .B(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hs__and2_2 _09021_ (.A(net2291),
    .B(net2298),
    .X(_03377_));
 sky130_fd_sc_hs__nand4_2 _09022_ (.A(_03372_),
    .B(_03374_),
    .C(_03376_),
    .D(net2281),
    .Y(_03378_));
 sky130_fd_sc_hs__xnor2_1 _09023_ (.A(_03344_),
    .B(net2331),
    .Y(_03379_));
 sky130_fd_sc_hs__nand2_1 _09024_ (.A(_03342_),
    .B(_03379_),
    .Y(_03380_));
 sky130_fd_sc_hs__nand3_1 _09025_ (.A(net2304),
    .B(net2331),
    .C(net2329),
    .Y(_03381_));
 sky130_fd_sc_hs__nand2_1 _09026_ (.A(_03380_),
    .B(_03381_),
    .Y(_03382_));
 sky130_fd_sc_hs__nand3b_1 _09027_ (.A_N(_03382_),
    .B(_03377_),
    .C(_03347_),
    .Y(_03383_));
 sky130_fd_sc_hs__nand2_2 _09028_ (.A(net2291),
    .B(net2298),
    .Y(_03384_));
 sky130_fd_sc_hs__o21ai_2 _09029_ (.A1(_03373_),
    .A2(_03384_),
    .B1(_03382_),
    .Y(_03385_));
 sky130_fd_sc_hs__nand2_1 _09030_ (.A(_03383_),
    .B(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hs__nand2_2 _09031_ (.A(_03371_),
    .B(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hs__nand3_2 _09032_ (.A(net5140),
    .B(_03370_),
    .C(net2280),
    .Y(_03388_));
 sky130_fd_sc_hs__nand2_2 _09033_ (.A(_03388_),
    .B(_03387_),
    .Y(_03389_));
 sky130_fd_sc_hs__o21ai_2 _09034_ (.A1(_03369_),
    .A2(_03365_),
    .B1(net2284),
    .Y(_03390_));
 sky130_fd_sc_hs__nand2_1 _09035_ (.A(_03390_),
    .B(net2282),
    .Y(_03391_));
 sky130_fd_sc_hs__and2b_1 _09036_ (.A_N(_03364_),
    .B(net5166),
    .X(_03392_));
 sky130_fd_sc_hs__nand2_2 _09037_ (.A(_03371_),
    .B(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hs__nand2_2 _09038_ (.A(_03391_),
    .B(_03393_),
    .Y(_03394_));
 sky130_fd_sc_hs__nor2_4 _09039_ (.A(_03394_),
    .B(_03389_),
    .Y(_03395_));
 sky130_fd_sc_hs__nand2_2 _09040_ (.A(_03378_),
    .B(_03395_),
    .Y(_03396_));
 sky130_fd_sc_hs__nand2_1 _09041_ (.A(_03393_),
    .B(net2283),
    .Y(_03397_));
 sky130_fd_sc_hs__nand2_1 _09042_ (.A(_03397_),
    .B(net2270),
    .Y(_03398_));
 sky130_fd_sc_hs__nand2_2 _09043_ (.A(_03396_),
    .B(_03398_),
    .Y(_03399_));
 sky130_fd_sc_hs__and2_1 _09044_ (.A(net2255),
    .B(net2265),
    .X(_03400_));
 sky130_fd_sc_hs__nand3_2 _09045_ (.A(_03399_),
    .B(_03376_),
    .C(_03400_),
    .Y(_03401_));
 sky130_fd_sc_hs__xnor2_1 _09046_ (.A(net2279),
    .B(net2255),
    .Y(_03402_));
 sky130_fd_sc_hs__nand2_1 _09047_ (.A(_03402_),
    .B(_03401_),
    .Y(_03403_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09048_ (.A(_03376_),
    .Y(_03404_));
 sky130_fd_sc_hs__nand3_1 _09049_ (.A(net2255),
    .B(net2264),
    .C(net2281),
    .Y(_03405_));
 sky130_fd_sc_hs__nor2_2 _09050_ (.A(_03404_),
    .B(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hs__nand2_1 _09051_ (.A(_03399_),
    .B(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hs__nand2_2 _09052_ (.A(_03407_),
    .B(_03403_),
    .Y(_03408_));
 sky130_fd_sc_hs__nand3_2 _09053_ (.A(_03396_),
    .B(_03376_),
    .C(_03398_),
    .Y(_03409_));
 sky130_fd_sc_hs__o21bai_1 _09054_ (.A1(net2282),
    .A2(net2269),
    .B1_N(net2283),
    .Y(_03410_));
 sky130_fd_sc_hs__nand3_1 _09055_ (.A(net2274),
    .B(net2290),
    .C(net2283),
    .Y(_03411_));
 sky130_fd_sc_hs__nand2_1 _09056_ (.A(_03410_),
    .B(_03411_),
    .Y(_03412_));
 sky130_fd_sc_hs__o21ai_2 _09057_ (.A1(_03412_),
    .A2(net2237),
    .B1(_03404_),
    .Y(_03413_));
 sky130_fd_sc_hs__nand2_2 _09058_ (.A(_03413_),
    .B(_03409_),
    .Y(_03414_));
 sky130_fd_sc_hs__nor2_1 _09059_ (.A(net3170),
    .B(net3132),
    .Y(_03415_));
 sky130_fd_sc_hs__xnor2_1 _09060_ (.A(net3260),
    .B(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09061_ (.A(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hs__nand3_2 _09062_ (.A(_03414_),
    .B(_03417_),
    .C(net2245),
    .Y(_03418_));
 sky130_fd_sc_hs__and2_1 _09063_ (.A(_03391_),
    .B(_03393_),
    .X(_03419_));
 sky130_fd_sc_hs__and2_1 _09064_ (.A(_03387_),
    .B(_03388_),
    .X(_03420_));
 sky130_fd_sc_hs__nand2_1 _09065_ (.A(_03419_),
    .B(_03420_),
    .Y(_03421_));
 sky130_fd_sc_hs__a21oi_1 _09066_ (.A1(_03421_),
    .A2(_03398_),
    .B1(_03406_),
    .Y(_03422_));
 sky130_fd_sc_hs__nand2_1 _09067_ (.A(_03422_),
    .B(net2247),
    .Y(_03423_));
 sky130_fd_sc_hs__o21ai_1 _09068_ (.A1(_03412_),
    .A2(net2236),
    .B1(net2248),
    .Y(_03424_));
 sky130_fd_sc_hs__nand2_1 _09069_ (.A(_03424_),
    .B(net2244),
    .Y(_03425_));
 sky130_fd_sc_hs__nand2_2 _09070_ (.A(_03423_),
    .B(_03425_),
    .Y(_03426_));
 sky130_fd_sc_hs__nand3_2 _09071_ (.A(_03418_),
    .B(_03426_),
    .C(_03408_),
    .Y(_03427_));
 sky130_fd_sc_hs__nand2_1 _09072_ (.A(net2248),
    .B(_03420_),
    .Y(_03428_));
 sky130_fd_sc_hs__o21ai_1 _09073_ (.A1(net2235),
    .A2(_03428_),
    .B1(net2246),
    .Y(_03429_));
 sky130_fd_sc_hs__and2_2 _09074_ (.A(_03429_),
    .B(net2231),
    .X(_03430_));
 sky130_fd_sc_hs__inv_4 _09075_ (.A(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hs__nand2_2 _09076_ (.A(_03427_),
    .B(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hs__xnor2_1 _09077_ (.A(_03416_),
    .B(net2215),
    .Y(_03433_));
 sky130_fd_sc_hs__nand2_1 _09078_ (.A(_03432_),
    .B(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hs__nand3_2 _09079_ (.A(net2194),
    .B(net2215),
    .C(net2213),
    .Y(_03435_));
 sky130_fd_sc_hs__nand2_2 _09080_ (.A(_03435_),
    .B(_03434_),
    .Y(_03436_));
 sky130_fd_sc_hs__nand2_1 _09081_ (.A(_03408_),
    .B(_03418_),
    .Y(_03437_));
 sky130_fd_sc_hs__inv_1 _09082_ (.A(net2214),
    .Y(_03438_));
 sky130_fd_sc_hs__o21ai_2 _09083_ (.A1(_03431_),
    .A2(_03437_),
    .B1(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hs__nand2_2 _09084_ (.A(_03439_),
    .B(net2194),
    .Y(_03440_));
 sky130_fd_sc_hs__and2_2 _09085_ (.A(_03436_),
    .B(_03440_),
    .X(_03441_));
 sky130_fd_sc_hs__o21ai_1 _09086_ (.A1(_02909_),
    .A2(net3334),
    .B1(net3089),
    .Y(_03442_));
 sky130_fd_sc_hs__xnor2_1 _09087_ (.A(net3333),
    .B(_03442_),
    .Y(_03443_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09088_ (.A(net2981),
    .Y(_03444_));
 sky130_fd_sc_hs__nand2_2 _09089_ (.A(_03432_),
    .B(_03417_),
    .Y(_03445_));
 sky130_fd_sc_hs__nand2_1 _09090_ (.A(_03408_),
    .B(_03426_),
    .Y(_03446_));
 sky130_fd_sc_hs__nand3_2 _09091_ (.A(_03446_),
    .B(_03416_),
    .C(_03431_),
    .Y(_03447_));
 sky130_fd_sc_hs__nand2_2 _09092_ (.A(_03445_),
    .B(_03447_),
    .Y(_03448_));
 sky130_fd_sc_hs__nor2_2 _09093_ (.A(_03444_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hs__nand2_2 _09094_ (.A(_03441_),
    .B(_03449_),
    .Y(_03450_));
 sky130_fd_sc_hs__o211ai_1 _09095_ (.A1(_03426_),
    .A2(_03430_),
    .B1(net2204),
    .C1(net5130),
    .Y(_03451_));
 sky130_fd_sc_hs__a21o_1 _09096_ (.A1(_03418_),
    .A2(_03430_),
    .B1(_03408_),
    .X(_03452_));
 sky130_fd_sc_hs__and2_2 _09097_ (.A(_03451_),
    .B(_03452_),
    .X(_03453_));
 sky130_fd_sc_hs__nand2_1 _09098_ (.A(net2226),
    .B(_03376_),
    .Y(_03454_));
 sky130_fd_sc_hs__inv_1 _09099_ (.A(net2245),
    .Y(_03455_));
 sky130_fd_sc_hs__nand2_1 _09100_ (.A(_03454_),
    .B(_03455_),
    .Y(_03456_));
 sky130_fd_sc_hs__nand2_1 _09101_ (.A(_03456_),
    .B(net2216),
    .Y(_03457_));
 sky130_fd_sc_hs__and2_1 _09102_ (.A(_03409_),
    .B(_03413_),
    .X(_03458_));
 sky130_fd_sc_hs__nor2_1 _09103_ (.A(_03416_),
    .B(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hs__xnor2_1 _09104_ (.A(_03457_),
    .B(_03459_),
    .Y(_03460_));
 sky130_fd_sc_hs__nand2_2 _09105_ (.A(_03432_),
    .B(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hs__inv_1 _09106_ (.A(net2198),
    .Y(_03462_));
 sky130_fd_sc_hs__nand3_1 _09107_ (.A(_03427_),
    .B(_03462_),
    .C(_03431_),
    .Y(_03463_));
 sky130_fd_sc_hs__nand3_1 _09108_ (.A(_03453_),
    .B(_03461_),
    .C(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hs__nand2_2 _09109_ (.A(_03464_),
    .B(_03440_),
    .Y(_03465_));
 sky130_fd_sc_hs__nand3_2 _09110_ (.A(_03450_),
    .B(_03444_),
    .C(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hs__nand2_1 _09111_ (.A(_03451_),
    .B(_03452_),
    .Y(_03467_));
 sky130_fd_sc_hs__nand2_2 _09112_ (.A(_03461_),
    .B(_03463_),
    .Y(_03468_));
 sky130_fd_sc_hs__nor2_2 _09113_ (.A(_03467_),
    .B(_03468_),
    .Y(_03469_));
 sky130_fd_sc_hs__nand3_1 _09114_ (.A(_03445_),
    .B(net2215),
    .C(_03447_),
    .Y(_03470_));
 sky130_fd_sc_hs__nand2_1 _09115_ (.A(_03469_),
    .B(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hs__nand3_2 _09116_ (.A(_03471_),
    .B(net2981),
    .C(net2177),
    .Y(_03472_));
 sky130_fd_sc_hs__nand2_2 _09117_ (.A(_03472_),
    .B(_03466_),
    .Y(_03473_));
 sky130_fd_sc_hs__or2_1 _09118_ (.A(net3167),
    .B(net3132),
    .X(_03474_));
 sky130_fd_sc_hs__xnor2_1 _09119_ (.A(net3294),
    .B(_03474_),
    .Y(_03475_));
 sky130_fd_sc_hs__inv_1 _09120_ (.A(net2163),
    .Y(_03476_));
 sky130_fd_sc_hs__nand3_2 _09121_ (.A(_03476_),
    .B(_03475_),
    .C(_03473_),
    .Y(_03477_));
 sky130_fd_sc_hs__nand4_2 _09122_ (.A(_03445_),
    .B(net2981),
    .C(net2215),
    .D(_03447_),
    .Y(_03478_));
 sky130_fd_sc_hs__and2_1 _09123_ (.A(_03439_),
    .B(net2194),
    .X(_03479_));
 sky130_fd_sc_hs__inv_1 _09124_ (.A(_03468_),
    .Y(_03480_));
 sky130_fd_sc_hs__a21o_1 _09125_ (.A1(_03478_),
    .A2(_03479_),
    .B1(_03480_),
    .X(_03481_));
 sky130_fd_sc_hs__o211ai_1 _09126_ (.A1(_03479_),
    .A2(net2187),
    .B1(_03480_),
    .C1(_03478_),
    .Y(_03482_));
 sky130_fd_sc_hs__nand2_2 _09127_ (.A(_03481_),
    .B(_03482_),
    .Y(_03483_));
 sky130_fd_sc_hs__nand3_1 _09128_ (.A(net5190),
    .B(net2981),
    .C(_03447_),
    .Y(_03484_));
 sky130_fd_sc_hs__nand2_1 _09129_ (.A(_03484_),
    .B(net2164),
    .Y(_03485_));
 sky130_fd_sc_hs__nand4_1 _09130_ (.A(_03445_),
    .B(net2981),
    .C(net2212),
    .D(net2188),
    .Y(_03486_));
 sky130_fd_sc_hs__nand2_1 _09131_ (.A(_03485_),
    .B(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hs__nand3_1 _09132_ (.A(_03487_),
    .B(_03450_),
    .C(net2156),
    .Y(_03488_));
 sky130_fd_sc_hs__nand2_2 _09133_ (.A(_03478_),
    .B(_03469_),
    .Y(_03489_));
 sky130_fd_sc_hs__nand3_1 _09134_ (.A(_03489_),
    .B(net2165),
    .C(net2177),
    .Y(_03490_));
 sky130_fd_sc_hs__nand2_2 _09135_ (.A(_03488_),
    .B(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hs__nor2_4 _09136_ (.A(_03483_),
    .B(_03491_),
    .Y(_03492_));
 sky130_fd_sc_hs__nand2_2 _09137_ (.A(_03492_),
    .B(_03477_),
    .Y(_03493_));
 sky130_fd_sc_hs__nand2_1 _09138_ (.A(_03482_),
    .B(net2186),
    .Y(_03494_));
 sky130_fd_sc_hs__nand2_2 _09139_ (.A(_03494_),
    .B(net2154),
    .Y(_03495_));
 sky130_fd_sc_hs__nand2_2 _09140_ (.A(_03493_),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09141_ (.A(_03475_),
    .Y(_03497_));
 sky130_fd_sc_hs__nand2_1 _09142_ (.A(_03473_),
    .B(_03476_),
    .Y(_03498_));
 sky130_fd_sc_hs__nor2_1 _09143_ (.A(_03497_),
    .B(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hs__nor2_1 _09144_ (.A(net2139),
    .B(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hs__nand2_2 _09145_ (.A(_03496_),
    .B(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hs__o21ai_1 _09146_ (.A1(_03495_),
    .A2(_03499_),
    .B1(net2139),
    .Y(_03502_));
 sky130_fd_sc_hs__and2_1 _09147_ (.A(_03501_),
    .B(_03502_),
    .X(_03503_));
 sky130_fd_sc_hs__inv_1 _09148_ (.A(net2139),
    .Y(_03504_));
 sky130_fd_sc_hs__nand2_1 _09149_ (.A(net2129),
    .B(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hs__o21ai_1 _09150_ (.A1(net2138),
    .A2(_03505_),
    .B1(net2146),
    .Y(_03506_));
 sky130_fd_sc_hs__and2_2 _09151_ (.A(_03506_),
    .B(net2122),
    .X(_03507_));
 sky130_fd_sc_hs__a21oi_1 _09152_ (.A1(net2157),
    .A2(net2981),
    .B1(_03476_),
    .Y(_03508_));
 sky130_fd_sc_hs__a21oi_4 _09153_ (.A1(net2154),
    .A2(net2177),
    .B1(net2162),
    .Y(_03509_));
 sky130_fd_sc_hs__nor2_2 _09154_ (.A(_03508_),
    .B(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hs__nand2_1 _09155_ (.A(net2140),
    .B(_03475_),
    .Y(_03511_));
 sky130_fd_sc_hs__xnor2_1 _09156_ (.A(_03510_),
    .B(_03511_),
    .Y(_03512_));
 sky130_fd_sc_hs__nand2_1 _09157_ (.A(_03512_),
    .B(_03496_),
    .Y(_03513_));
 sky130_fd_sc_hs__nand3_1 _09158_ (.A(_03493_),
    .B(_03510_),
    .C(_03495_),
    .Y(_03514_));
 sky130_fd_sc_hs__nand2_2 _09159_ (.A(_03513_),
    .B(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hs__inv_1 _09160_ (.A(net2104),
    .Y(_03516_));
 sky130_fd_sc_hs__nand2_2 _09161_ (.A(_03496_),
    .B(_03475_),
    .Y(_03517_));
 sky130_fd_sc_hs__nand3_2 _09162_ (.A(net5120),
    .B(_03497_),
    .C(net2137),
    .Y(_03518_));
 sky130_fd_sc_hs__nor2_1 _09163_ (.A(net3262),
    .B(net3132),
    .Y(_03519_));
 sky130_fd_sc_hs__xnor2_1 _09164_ (.A(net3382),
    .B(_03519_),
    .Y(_03520_));
 sky130_fd_sc_hs__nand4_2 _09165_ (.A(_03517_),
    .B(_03518_),
    .C(_03520_),
    .D(net2140),
    .Y(_03521_));
 sky130_fd_sc_hs__o211ai_1 _09166_ (.A1(_03503_),
    .A2(_03507_),
    .B1(_03516_),
    .C1(net2103),
    .Y(_03522_));
 sky130_fd_sc_hs__nand2_2 _09167_ (.A(_03501_),
    .B(_03502_),
    .Y(_03523_));
 sky130_fd_sc_hs__nand2_1 _09168_ (.A(_03522_),
    .B(net2102),
    .Y(_03524_));
 sky130_fd_sc_hs__nor2_4 _09169_ (.A(_03515_),
    .B(_03523_),
    .Y(_03525_));
 sky130_fd_sc_hs__nand2_2 _09170_ (.A(_03521_),
    .B(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hs__nand2_4 _09171_ (.A(_03524_),
    .B(net2087),
    .Y(_03527_));
 sky130_fd_sc_hs__inv_1 _09172_ (.A(_03507_),
    .Y(_03528_));
 sky130_fd_sc_hs__nand2_2 _09173_ (.A(_03528_),
    .B(_03526_),
    .Y(_03529_));
 sky130_fd_sc_hs__nand2_2 _09174_ (.A(_03529_),
    .B(_03520_),
    .Y(_03530_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09175_ (.A(_03520_),
    .Y(_03531_));
 sky130_fd_sc_hs__nand3_2 _09176_ (.A(_03526_),
    .B(_03531_),
    .C(_03528_),
    .Y(_03532_));
 sky130_fd_sc_hs__and2_1 _09177_ (.A(net3090),
    .B(net3381),
    .X(_03533_));
 sky130_fd_sc_hs__xnor2_1 _09178_ (.A(net3295),
    .B(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09179_ (.A(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hs__nand2_1 _09180_ (.A(net2111),
    .B(net2119),
    .Y(_03536_));
 sky130_fd_sc_hs__nor2_1 _09181_ (.A(_03535_),
    .B(_03536_),
    .Y(_03537_));
 sky130_fd_sc_hs__nand3_4 _09182_ (.A(_03532_),
    .B(_03530_),
    .C(_03537_),
    .Y(_03538_));
 sky130_fd_sc_hs__xnor2_1 _09183_ (.A(_03497_),
    .B(net2140),
    .Y(_03539_));
 sky130_fd_sc_hs__nand2_1 _09184_ (.A(_03496_),
    .B(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hs__nand3_1 _09185_ (.A(_03493_),
    .B(net2140),
    .C(_03495_),
    .Y(_03541_));
 sky130_fd_sc_hs__nand2_1 _09186_ (.A(_03540_),
    .B(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hs__nand3_2 _09187_ (.A(net2111),
    .B(net2119),
    .C(_03520_),
    .Y(_03543_));
 sky130_fd_sc_hs__xnor2_2 _09188_ (.A(_03543_),
    .B(_03542_),
    .Y(_03544_));
 sky130_fd_sc_hs__nand2_1 _09189_ (.A(_03544_),
    .B(_03529_),
    .Y(_03545_));
 sky130_fd_sc_hs__nand3_1 _09190_ (.A(_03526_),
    .B(_03528_),
    .C(net2100),
    .Y(_03546_));
 sky130_fd_sc_hs__and2_1 _09191_ (.A(_03545_),
    .B(_03546_),
    .X(_03547_));
 sky130_fd_sc_hs__nand2_2 _09192_ (.A(_03538_),
    .B(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hs__a21o_1 _09193_ (.A1(net2103),
    .A2(_03507_),
    .B1(_03516_),
    .X(_03549_));
 sky130_fd_sc_hs__nand2_1 _09194_ (.A(_03522_),
    .B(_03549_),
    .Y(_03550_));
 sky130_fd_sc_hs__o21ai_1 _09195_ (.A1(_03527_),
    .A2(_03548_),
    .B1(net2081),
    .Y(_03551_));
 sky130_fd_sc_hs__nand2_1 _09196_ (.A(_03545_),
    .B(_03546_),
    .Y(_03552_));
 sky130_fd_sc_hs__nor2_2 _09197_ (.A(_03550_),
    .B(_03552_),
    .Y(_03553_));
 sky130_fd_sc_hs__nand2_2 _09198_ (.A(_03538_),
    .B(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hs__and2_2 _09199_ (.A(_03551_),
    .B(net5131),
    .X(_03555_));
 sky130_fd_sc_hs__a21o_1 _09200_ (.A1(_03527_),
    .A2(net2081),
    .B1(_03548_),
    .X(_03556_));
 sky130_fd_sc_hs__and2_1 _09201_ (.A(_03524_),
    .B(net2087),
    .X(_03557_));
 sky130_fd_sc_hs__a21o_1 _09202_ (.A1(_03557_),
    .A2(_03538_),
    .B1(_03547_),
    .X(_03558_));
 sky130_fd_sc_hs__and2_1 _09203_ (.A(_03556_),
    .B(_03558_),
    .X(_03559_));
 sky130_fd_sc_hs__nand2_1 _09204_ (.A(_03530_),
    .B(net2082),
    .Y(_03560_));
 sky130_fd_sc_hs__xnor2_1 _09205_ (.A(_03520_),
    .B(_03536_),
    .Y(_03561_));
 sky130_fd_sc_hs__nand2_1 _09206_ (.A(net2085),
    .B(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hs__o21ai_2 _09207_ (.A1(_03536_),
    .A2(net2084),
    .B1(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hs__o21ai_1 _09208_ (.A1(_03535_),
    .A2(_03560_),
    .B1(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hs__nand4_1 _09209_ (.A(net2072),
    .B(net2082),
    .C(_03534_),
    .D(net2101),
    .Y(_03565_));
 sky130_fd_sc_hs__nand2_1 _09210_ (.A(_03564_),
    .B(_03565_),
    .Y(_03566_));
 sky130_fd_sc_hs__nand2_2 _09211_ (.A(_03554_),
    .B(_03527_),
    .Y(_03567_));
 sky130_fd_sc_hs__nand2_2 _09212_ (.A(_03566_),
    .B(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hs__nand3_1 _09213_ (.A(_03554_),
    .B(net2073),
    .C(net2065),
    .Y(_03569_));
 sky130_fd_sc_hs__nand2_2 _09214_ (.A(_03568_),
    .B(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hs__inv_1 _09215_ (.A(_03570_),
    .Y(_03571_));
 sky130_fd_sc_hs__nand2_2 _09216_ (.A(_03567_),
    .B(_03534_),
    .Y(_03572_));
 sky130_fd_sc_hs__nand3_2 _09217_ (.A(_03554_),
    .B(_03535_),
    .C(_03527_),
    .Y(_03573_));
 sky130_fd_sc_hs__and2_1 _09218_ (.A(net3090),
    .B(net3443),
    .X(_03574_));
 sky130_fd_sc_hs__xnor2_1 _09219_ (.A(net3501),
    .B(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hs__and2_1 _09220_ (.A(net2072),
    .B(net2083),
    .X(_03576_));
 sky130_fd_sc_hs__nand4_2 _09221_ (.A(_03572_),
    .B(_03573_),
    .C(_03575_),
    .D(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hs__o211ai_2 _09222_ (.A1(_03555_),
    .A2(_03559_),
    .B1(_03571_),
    .C1(net2023),
    .Y(_03578_));
 sky130_fd_sc_hs__nand2_1 _09223_ (.A(_03556_),
    .B(_03558_),
    .Y(_03579_));
 sky130_fd_sc_hs__nand2_1 _09224_ (.A(_03578_),
    .B(net2046),
    .Y(_03580_));
 sky130_fd_sc_hs__nor2_4 _09225_ (.A(_03579_),
    .B(_03570_),
    .Y(_03581_));
 sky130_fd_sc_hs__nand2_2 _09226_ (.A(_03581_),
    .B(_03577_),
    .Y(_03582_));
 sky130_fd_sc_hs__nand2_4 _09227_ (.A(_03580_),
    .B(net2004),
    .Y(_03583_));
 sky130_fd_sc_hs__inv_8 _09228_ (.A(_03555_),
    .Y(_03584_));
 sky130_fd_sc_hs__nand2_2 _09229_ (.A(_03582_),
    .B(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hs__nand2_2 _09230_ (.A(_03585_),
    .B(_03575_),
    .Y(_03586_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09231_ (.A(_03575_),
    .Y(_03587_));
 sky130_fd_sc_hs__nand3_2 _09232_ (.A(net5126),
    .B(_03587_),
    .C(_03584_),
    .Y(_03588_));
 sky130_fd_sc_hs__nand2_1 _09233_ (.A(net3090),
    .B(net3380),
    .Y(_03589_));
 sky130_fd_sc_hs__xnor2_1 _09234_ (.A(net5174),
    .B(_03589_),
    .Y(_03590_));
 sky130_fd_sc_hs__nand2_1 _09235_ (.A(_03572_),
    .B(net2047),
    .Y(_03591_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09236_ (.A(_03591_),
    .Y(_03592_));
 sky130_fd_sc_hs__nand4_2 _09237_ (.A(_03586_),
    .B(_03588_),
    .C(_03590_),
    .D(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hs__nand2_1 _09238_ (.A(net2036),
    .B(net2066),
    .Y(_03594_));
 sky130_fd_sc_hs__nand3_1 _09239_ (.A(_03567_),
    .B(_03534_),
    .C(_03576_),
    .Y(_03595_));
 sky130_fd_sc_hs__nand2_2 _09240_ (.A(_03594_),
    .B(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hs__nor2_2 _09241_ (.A(_03587_),
    .B(_03591_),
    .Y(_03597_));
 sky130_fd_sc_hs__xnor2_1 _09242_ (.A(_03596_),
    .B(_03597_),
    .Y(_03598_));
 sky130_fd_sc_hs__nand2_1 _09243_ (.A(_03598_),
    .B(_03585_),
    .Y(_03599_));
 sky130_fd_sc_hs__nand3b_1 _09244_ (.A_N(net2011),
    .B(_03582_),
    .C(_03584_),
    .Y(_03600_));
 sky130_fd_sc_hs__nand2_2 _09245_ (.A(_03599_),
    .B(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hs__clkinv_1 _09246_ (.A(_03601_),
    .Y(_03602_));
 sky130_fd_sc_hs__nand2_1 _09247_ (.A(net5119),
    .B(_03602_),
    .Y(_03603_));
 sky130_fd_sc_hs__o21ai_1 _09248_ (.A1(_03555_),
    .A2(_03581_),
    .B1(net2023),
    .Y(_03604_));
 sky130_fd_sc_hs__nand2_1 _09249_ (.A(_03604_),
    .B(net2024),
    .Y(_03605_));
 sky130_fd_sc_hs__nand2_2 _09250_ (.A(_03578_),
    .B(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hs__o21ai_1 _09251_ (.A1(_03583_),
    .A2(_03603_),
    .B1(net1987),
    .Y(_03607_));
 sky130_fd_sc_hs__nor2_2 _09252_ (.A(_03606_),
    .B(_03601_),
    .Y(_03608_));
 sky130_fd_sc_hs__nand2_2 _09253_ (.A(_03608_),
    .B(_03593_),
    .Y(_03609_));
 sky130_fd_sc_hs__and2_1 _09254_ (.A(_03607_),
    .B(_03609_),
    .X(_03610_));
 sky130_fd_sc_hs__and2_1 _09255_ (.A(_03605_),
    .B(_03578_),
    .X(_03611_));
 sky130_fd_sc_hs__and2_1 _09256_ (.A(_03580_),
    .B(net2004),
    .X(_03612_));
 sky130_fd_sc_hs__o211ai_1 _09257_ (.A1(_03611_),
    .A2(_03612_),
    .B1(_03602_),
    .C1(net1981),
    .Y(_03613_));
 sky130_fd_sc_hs__a21o_1 _09258_ (.A1(net5119),
    .A2(_03612_),
    .B1(_03602_),
    .X(_03614_));
 sky130_fd_sc_hs__nand2_4 _09259_ (.A(_03613_),
    .B(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hs__nand2_2 _09260_ (.A(_03583_),
    .B(_03609_),
    .Y(_03616_));
 sky130_fd_sc_hs__nand2_1 _09261_ (.A(net1988),
    .B(net2022),
    .Y(_03617_));
 sky130_fd_sc_hs__nand2_1 _09262_ (.A(_03585_),
    .B(net2010),
    .Y(_03618_));
 sky130_fd_sc_hs__and2_2 _09263_ (.A(_03617_),
    .B(_03618_),
    .X(_03619_));
 sky130_fd_sc_hs__and2_2 _09264_ (.A(net1999),
    .B(net1988),
    .X(_03620_));
 sky130_fd_sc_hs__nand2_1 _09265_ (.A(_03620_),
    .B(_03590_),
    .Y(_03621_));
 sky130_fd_sc_hs__nand2_1 _09266_ (.A(_03621_),
    .B(_03619_),
    .Y(_03622_));
 sky130_fd_sc_hs__nand4_1 _09267_ (.A(net1989),
    .B(net1999),
    .C(_03590_),
    .D(net2022),
    .Y(_03623_));
 sky130_fd_sc_hs__nand2_1 _09268_ (.A(_03622_),
    .B(_03623_),
    .Y(_03624_));
 sky130_fd_sc_hs__nand2_2 _09269_ (.A(_03616_),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hs__nand3_1 _09270_ (.A(_03609_),
    .B(_03619_),
    .C(_03583_),
    .Y(_03626_));
 sky130_fd_sc_hs__nand2_2 _09271_ (.A(_03625_),
    .B(_03626_),
    .Y(_03627_));
 sky130_fd_sc_hs__nor2_4 _09272_ (.A(_03627_),
    .B(_03615_),
    .Y(_03628_));
 sky130_fd_sc_hs__nand2_2 _09273_ (.A(_03616_),
    .B(_03590_),
    .Y(_03629_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09274_ (.A(_03590_),
    .Y(_03630_));
 sky130_fd_sc_hs__nand3_2 _09275_ (.A(_03609_),
    .B(_03630_),
    .C(_03583_),
    .Y(_03631_));
 sky130_fd_sc_hs__o31ai_1 _09276_ (.A1(net3765),
    .A2(net3751),
    .A3(net3754),
    .B1(net3090),
    .Y(_03632_));
 sky130_fd_sc_hs__xnor2_1 _09277_ (.A(net3750),
    .B(_03632_),
    .Y(_03633_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09278_ (.A(_03633_),
    .Y(_03634_));
 sky130_fd_sc_hs__nand4_4 _09279_ (.A(_03629_),
    .B(_03631_),
    .C(_03634_),
    .D(net1980),
    .Y(_03635_));
 sky130_fd_sc_hs__o21ai_1 _09280_ (.A1(_03610_),
    .A2(net1926),
    .B1(net1938),
    .Y(_03636_));
 sky130_fd_sc_hs__inv_1 _09281_ (.A(net1939),
    .Y(_03637_));
 sky130_fd_sc_hs__nand2_1 _09282_ (.A(_03637_),
    .B(_03636_),
    .Y(_03638_));
 sky130_fd_sc_hs__nand3_1 _09283_ (.A(net1938),
    .B(net1939),
    .C(net1948),
    .Y(_03639_));
 sky130_fd_sc_hs__nand2_1 _09284_ (.A(_03639_),
    .B(_03638_),
    .Y(_03640_));
 sky130_fd_sc_hs__nand2_2 _09285_ (.A(_03635_),
    .B(_03628_),
    .Y(_03641_));
 sky130_fd_sc_hs__inv_4 _09286_ (.A(_03610_),
    .Y(_03642_));
 sky130_fd_sc_hs__nand2_2 _09287_ (.A(_03642_),
    .B(_03641_),
    .Y(_03643_));
 sky130_fd_sc_hs__nand2_1 _09288_ (.A(net1989),
    .B(net1999),
    .Y(_03644_));
 sky130_fd_sc_hs__nand2_1 _09289_ (.A(_03629_),
    .B(_03644_),
    .Y(_03645_));
 sky130_fd_sc_hs__nor2_1 _09290_ (.A(_03630_),
    .B(_03644_),
    .Y(_03646_));
 sky130_fd_sc_hs__nand2_1 _09291_ (.A(net1958),
    .B(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hs__and2_2 _09292_ (.A(_03645_),
    .B(_03647_),
    .X(_03648_));
 sky130_fd_sc_hs__nand3_1 _09293_ (.A(_03629_),
    .B(net1957),
    .C(_03634_),
    .Y(_03649_));
 sky130_fd_sc_hs__nand2_1 _09294_ (.A(_03648_),
    .B(_03649_),
    .Y(_03650_));
 sky130_fd_sc_hs__nand4_1 _09295_ (.A(_03629_),
    .B(net1957),
    .C(_03634_),
    .D(net1979),
    .Y(_03651_));
 sky130_fd_sc_hs__nand2_4 _09296_ (.A(_03650_),
    .B(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hs__nand2_2 _09297_ (.A(_03643_),
    .B(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hs__nand3_1 _09298_ (.A(_03641_),
    .B(net1925),
    .C(_03642_),
    .Y(_03654_));
 sky130_fd_sc_hs__nand2_2 _09299_ (.A(_03654_),
    .B(_03653_),
    .Y(_03655_));
 sky130_fd_sc_hs__and2b_2 _09300_ (.A_N(_03640_),
    .B(_03655_),
    .X(_03656_));
 sky130_fd_sc_hs__nand2_2 _09301_ (.A(_03643_),
    .B(_03634_),
    .Y(_03657_));
 sky130_fd_sc_hs__nand3_2 _09302_ (.A(_03642_),
    .B(_03633_),
    .C(_03641_),
    .Y(_03658_));
 sky130_fd_sc_hs__inv_1 _09303_ (.A(net3751),
    .Y(_03659_));
 sky130_fd_sc_hs__nor2_1 _09304_ (.A(net3421),
    .B(net3132),
    .Y(_03660_));
 sky130_fd_sc_hs__xnor2_1 _09305_ (.A(_03659_),
    .B(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09306_ (.A(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hs__nand3_1 _09307_ (.A(_03662_),
    .B(net3608),
    .C(_00215_),
    .Y(_03663_));
 sky130_fd_sc_hs__nand2_1 _09308_ (.A(_03629_),
    .B(net1957),
    .Y(_03664_));
 sky130_fd_sc_hs__nor2_1 _09309_ (.A(_03663_),
    .B(net1937),
    .Y(_03665_));
 sky130_fd_sc_hs__and3_4 _09310_ (.A(_03657_),
    .B(net5135),
    .C(_03665_),
    .X(_03666_));
 sky130_fd_sc_hs__a21o_1 _09311_ (.A1(net1938),
    .A2(_03637_),
    .B1(net1959),
    .X(_03667_));
 sky130_fd_sc_hs__nand4_1 _09312_ (.A(net1938),
    .B(_03637_),
    .C(net1959),
    .D(net1948),
    .Y(_03668_));
 sky130_fd_sc_hs__nand2_1 _09313_ (.A(_03667_),
    .B(_03668_),
    .Y(_03669_));
 sky130_fd_sc_hs__inv_4 _09314_ (.A(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hs__nand3_2 _09315_ (.A(_03656_),
    .B(_03666_),
    .C(_03670_),
    .Y(_03671_));
 sky130_fd_sc_hs__buf_1 place2129 (.A(_03477_),
    .X(net2129));
 sky130_fd_sc_hs__nand3_2 _09317_ (.A(net3777),
    .B(_03671_),
    .C(net3090),
    .Y(_03673_));
 sky130_fd_sc_hs__buf_1 place2128 (.A(_04575_),
    .X(net2128));
 sky130_fd_sc_hs__buf_1 place2126 (.A(_04588_),
    .X(net2126));
 sky130_fd_sc_hs__nand2_1 _09320_ (.A(net3673),
    .B(net3776),
    .Y(_03676_));
 sky130_fd_sc_hs__a21oi_2 _09321_ (.A1(net1874),
    .A2(_03676_),
    .B1(net3783),
    .Y(_00428_));
 sky130_fd_sc_hs__and2_1 _09322_ (.A(_03638_),
    .B(_03639_),
    .X(_03677_));
 sky130_fd_sc_hs__nand2_1 _09323_ (.A(_03670_),
    .B(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hs__xnor2_1 _09324_ (.A(_03634_),
    .B(_03664_),
    .Y(_03679_));
 sky130_fd_sc_hs__nand2_1 _09325_ (.A(_03643_),
    .B(_03679_),
    .Y(_03680_));
 sky130_fd_sc_hs__inv_1 _09326_ (.A(_03664_),
    .Y(_03681_));
 sky130_fd_sc_hs__nand3_1 _09327_ (.A(_03641_),
    .B(_03681_),
    .C(_03642_),
    .Y(_03682_));
 sky130_fd_sc_hs__nand2_2 _09328_ (.A(_03680_),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hs__and2_2 _09329_ (.A(_03655_),
    .B(_03683_),
    .X(_03684_));
 sky130_fd_sc_hs__and2_1 _09330_ (.A(_03662_),
    .B(_00216_),
    .X(_03685_));
 sky130_fd_sc_hs__and3_2 _09331_ (.A(_03658_),
    .B(_03657_),
    .C(_03685_),
    .X(_03686_));
 sky130_fd_sc_hs__nand2_2 _09332_ (.A(_03686_),
    .B(_03684_),
    .Y(_03687_));
 sky130_fd_sc_hs__o211ai_4 _09333_ (.A1(_03678_),
    .A2(_03687_),
    .B1(net3777),
    .C1(net3090),
    .Y(_03688_));
 sky130_fd_sc_hs__buf_1 place2125 (.A(_05485_),
    .X(net2125));
 sky130_fd_sc_hs__nand2_1 _09335_ (.A(net3673),
    .B(net3775),
    .Y(_03690_));
 sky130_fd_sc_hs__a21oi_2 _09336_ (.A1(net1873),
    .A2(_03690_),
    .B1(net3783),
    .Y(_00429_));
 sky130_fd_sc_hs__nand2_1 _09337_ (.A(net3673),
    .B(net3774),
    .Y(_03691_));
 sky130_fd_sc_hs__buf_1 place2122 (.A(net5118),
    .X(net2122));
 sky130_fd_sc_hs__a21oi_2 _09339_ (.A1(net1874),
    .A2(_03691_),
    .B1(net3783),
    .Y(_00430_));
 sky130_fd_sc_hs__nand2_1 _09340_ (.A(net3673),
    .B(net3773),
    .Y(_03693_));
 sky130_fd_sc_hs__a21oi_2 _09341_ (.A1(net1873),
    .A2(_03693_),
    .B1(net3783),
    .Y(_00431_));
 sky130_fd_sc_hs__nand2_1 _09342_ (.A(net3673),
    .B(net3771),
    .Y(_03694_));
 sky130_fd_sc_hs__a21oi_2 _09343_ (.A1(net1874),
    .A2(_03694_),
    .B1(net3783),
    .Y(_00432_));
 sky130_fd_sc_hs__nand2_1 _09344_ (.A(net3673),
    .B(net3770),
    .Y(_03695_));
 sky130_fd_sc_hs__a21oi_2 _09345_ (.A1(net1873),
    .A2(_03695_),
    .B1(net3783),
    .Y(_00433_));
 sky130_fd_sc_hs__nand2_1 _09346_ (.A(net3673),
    .B(net3769),
    .Y(_03696_));
 sky130_fd_sc_hs__a21oi_2 _09347_ (.A1(net1874),
    .A2(_03696_),
    .B1(net3783),
    .Y(_00434_));
 sky130_fd_sc_hs__nand2_1 _09348_ (.A(net3673),
    .B(net3768),
    .Y(_03697_));
 sky130_fd_sc_hs__a21oi_2 _09349_ (.A1(net1873),
    .A2(_03697_),
    .B1(net3783),
    .Y(_00435_));
 sky130_fd_sc_hs__buf_1 place2121 (.A(net5095),
    .X(net2121));
 sky130_fd_sc_hs__nand2_1 _09351_ (.A(net3673),
    .B(net3767),
    .Y(_03699_));
 sky130_fd_sc_hs__a21oi_2 _09352_ (.A1(net1874),
    .A2(_03699_),
    .B1(net3783),
    .Y(_00436_));
 sky130_fd_sc_hs__nand2_1 _09353_ (.A(net3673),
    .B(net3766),
    .Y(_03700_));
 sky130_fd_sc_hs__a21oi_2 _09354_ (.A1(net1873),
    .A2(_03700_),
    .B1(net3783),
    .Y(_00437_));
 sky130_fd_sc_hs__o21ai_1 _09355_ (.A1(\u_window_buffer.current_state[3] ),
    .A2(_00658_),
    .B1(net3765),
    .Y(_03701_));
 sky130_fd_sc_hs__nor2_1 _09356_ (.A(net3782),
    .B(_03701_),
    .Y(_00438_));
 sky130_fd_sc_hs__nand2_1 _09357_ (.A(net3673),
    .B(net3764),
    .Y(_03702_));
 sky130_fd_sc_hs__a21oi_2 _09358_ (.A1(net1874),
    .A2(_03702_),
    .B1(net3783),
    .Y(_00439_));
 sky130_fd_sc_hs__nand2_1 _09359_ (.A(net3673),
    .B(net3763),
    .Y(_03703_));
 sky130_fd_sc_hs__a21oi_2 _09360_ (.A1(net1873),
    .A2(_03703_),
    .B1(net3783),
    .Y(_00440_));
 sky130_fd_sc_hs__nand2_1 _09361_ (.A(net3673),
    .B(net3762),
    .Y(_03704_));
 sky130_fd_sc_hs__buf_1 place2120 (.A(_01740_),
    .X(net2120));
 sky130_fd_sc_hs__a21oi_2 _09363_ (.A1(net1874),
    .A2(_03704_),
    .B1(net3783),
    .Y(_00441_));
 sky130_fd_sc_hs__nand2_1 _09364_ (.A(net3673),
    .B(net3761),
    .Y(_03706_));
 sky130_fd_sc_hs__a21oi_2 _09365_ (.A1(net1873),
    .A2(_03706_),
    .B1(net3783),
    .Y(_00442_));
 sky130_fd_sc_hs__nand2_1 _09366_ (.A(net3673),
    .B(net3760),
    .Y(_03707_));
 sky130_fd_sc_hs__a21oi_2 _09367_ (.A1(net1874),
    .A2(_03707_),
    .B1(net3783),
    .Y(_00443_));
 sky130_fd_sc_hs__nand2_1 _09368_ (.A(net3673),
    .B(net3759),
    .Y(_03708_));
 sky130_fd_sc_hs__a21oi_2 _09369_ (.A1(net1873),
    .A2(_03708_),
    .B1(net3783),
    .Y(_00444_));
 sky130_fd_sc_hs__nand2_1 _09370_ (.A(net3673),
    .B(net3758),
    .Y(_03709_));
 sky130_fd_sc_hs__a21oi_2 _09371_ (.A1(net1874),
    .A2(_03709_),
    .B1(net3783),
    .Y(_00445_));
 sky130_fd_sc_hs__nand2_1 _09372_ (.A(net3673),
    .B(net3757),
    .Y(_03710_));
 sky130_fd_sc_hs__a21oi_2 _09373_ (.A1(net1873),
    .A2(_03710_),
    .B1(net3783),
    .Y(_00446_));
 sky130_fd_sc_hs__buf_1 place2119 (.A(_03518_),
    .X(net2119));
 sky130_fd_sc_hs__nand2_1 _09375_ (.A(net3673),
    .B(net3756),
    .Y(_03712_));
 sky130_fd_sc_hs__a21oi_2 _09376_ (.A1(net1874),
    .A2(_03712_),
    .B1(net3783),
    .Y(_00447_));
 sky130_fd_sc_hs__nand2_1 _09377_ (.A(net3673),
    .B(net3755),
    .Y(_03713_));
 sky130_fd_sc_hs__a21oi_2 _09378_ (.A1(net1873),
    .A2(_03713_),
    .B1(net3783),
    .Y(_00448_));
 sky130_fd_sc_hs__o21ai_1 _09379_ (.A1(_00217_),
    .A2(net3132),
    .B1(net3777),
    .Y(_03714_));
 sky130_fd_sc_hs__nand2_1 _09380_ (.A(net3673),
    .B(net3754),
    .Y(_03715_));
 sky130_fd_sc_hs__a211oi_1 _09381_ (.A1(_03714_),
    .A2(_03715_),
    .B1(net3783),
    .C1(_02235_),
    .Y(_00449_));
 sky130_fd_sc_hs__nand2_1 _09382_ (.A(net3673),
    .B(net3753),
    .Y(_03716_));
 sky130_fd_sc_hs__a21oi_1 _09383_ (.A1(net1874),
    .A2(_03716_),
    .B1(net3783),
    .Y(_00450_));
 sky130_fd_sc_hs__nand2_1 _09384_ (.A(net3673),
    .B(net3752),
    .Y(_03717_));
 sky130_fd_sc_hs__a21oi_1 _09385_ (.A1(net1873),
    .A2(_03717_),
    .B1(net3783),
    .Y(_00451_));
 sky130_fd_sc_hs__nor2_1 _09386_ (.A(_00216_),
    .B(_03662_),
    .Y(_03718_));
 sky130_fd_sc_hs__o21ai_1 _09387_ (.A1(_03718_),
    .A2(_03685_),
    .B1(net3090),
    .Y(_03719_));
 sky130_fd_sc_hs__o211ai_1 _09388_ (.A1(net3751),
    .A2(net3090),
    .B1(net3777),
    .C1(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hs__nand2_1 _09389_ (.A(net3673),
    .B(net3751),
    .Y(_03721_));
 sky130_fd_sc_hs__a21oi_1 _09390_ (.A1(_03720_),
    .A2(_03721_),
    .B1(net3783),
    .Y(_00452_));
 sky130_fd_sc_hs__nand2_1 _09391_ (.A(net1912),
    .B(net1921),
    .Y(_03722_));
 sky130_fd_sc_hs__and2_1 _09392_ (.A(_03663_),
    .B(net3090),
    .X(_03723_));
 sky130_fd_sc_hs__o21ai_1 _09393_ (.A1(_03723_),
    .A2(_03722_),
    .B1(net3777),
    .Y(_03724_));
 sky130_fd_sc_hs__a21o_1 _09394_ (.A1(_03722_),
    .A2(_03723_),
    .B1(_03724_),
    .X(_03725_));
 sky130_fd_sc_hs__nand2_1 _09395_ (.A(net3673),
    .B(net3750),
    .Y(_03726_));
 sky130_fd_sc_hs__a21oi_4 _09396_ (.A1(_03726_),
    .A2(_03725_),
    .B1(net3783),
    .Y(_00453_));
 sky130_fd_sc_hs__nor3_2 _09397_ (.A(net3132),
    .B(net1900),
    .C(net5262),
    .Y(_03727_));
 sky130_fd_sc_hs__o21ai_2 _09398_ (.A1(net3132),
    .A2(net5262),
    .B1(net1900),
    .Y(_03728_));
 sky130_fd_sc_hs__nand3b_1 _09399_ (.A_N(_03727_),
    .B(net3777),
    .C(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hs__nand2_1 _09400_ (.A(net3673),
    .B(net3749),
    .Y(_03730_));
 sky130_fd_sc_hs__a21oi_1 _09401_ (.A1(_03730_),
    .A2(_03729_),
    .B1(net3783),
    .Y(_00454_));
 sky130_fd_sc_hs__nor3_2 _09402_ (.A(net3132),
    .B(_03666_),
    .C(net1901),
    .Y(_03731_));
 sky130_fd_sc_hs__o21ai_2 _09403_ (.A1(net3132),
    .A2(_03666_),
    .B1(net1901),
    .Y(_03732_));
 sky130_fd_sc_hs__nand3b_2 _09404_ (.A_N(_03731_),
    .B(net3777),
    .C(_03732_),
    .Y(_03733_));
 sky130_fd_sc_hs__nand2_1 _09405_ (.A(net3673),
    .B(net3748),
    .Y(_03734_));
 sky130_fd_sc_hs__a21oi_4 _09406_ (.A1(_03734_),
    .A2(_03733_),
    .B1(net3783),
    .Y(_00455_));
 sky130_fd_sc_hs__nand3_1 _09407_ (.A(_03657_),
    .B(net1920),
    .C(_03685_),
    .Y(_03735_));
 sky130_fd_sc_hs__nand2_1 _09408_ (.A(_03655_),
    .B(_03683_),
    .Y(_03736_));
 sky130_fd_sc_hs__o21ai_1 _09409_ (.A1(_03735_),
    .A2(_03736_),
    .B1(net3090),
    .Y(_03737_));
 sky130_fd_sc_hs__nand2_1 _09410_ (.A(_03737_),
    .B(net1909),
    .Y(_03738_));
 sky130_fd_sc_hs__nand3_1 _09411_ (.A(_03687_),
    .B(net3090),
    .C(net1913),
    .Y(_03739_));
 sky130_fd_sc_hs__nand3_2 _09412_ (.A(_03739_),
    .B(_03738_),
    .C(net3777),
    .Y(_03740_));
 sky130_fd_sc_hs__nand2_1 _09413_ (.A(net3673),
    .B(net3747),
    .Y(_03741_));
 sky130_fd_sc_hs__a21oi_4 _09414_ (.A1(_03741_),
    .A2(_03740_),
    .B1(net3783),
    .Y(_00456_));
 sky130_fd_sc_hs__nand3_2 _09415_ (.A(net1911),
    .B(net1919),
    .C(net1924),
    .Y(_03742_));
 sky130_fd_sc_hs__nand2_1 _09416_ (.A(_03677_),
    .B(_03655_),
    .Y(_03743_));
 sky130_fd_sc_hs__o21ai_2 _09417_ (.A1(_03743_),
    .A2(_03742_),
    .B1(net3090),
    .Y(_03744_));
 sky130_fd_sc_hs__nand2_1 _09418_ (.A(net1910),
    .B(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hs__nand2_1 _09419_ (.A(_03656_),
    .B(_03666_),
    .Y(_03746_));
 sky130_fd_sc_hs__nand3_1 _09420_ (.A(_03746_),
    .B(net3090),
    .C(net1918),
    .Y(_03747_));
 sky130_fd_sc_hs__nand3_2 _09421_ (.A(_03747_),
    .B(_03745_),
    .C(net3777),
    .Y(_03748_));
 sky130_fd_sc_hs__nand2_1 _09422_ (.A(_00658_),
    .B(net3746),
    .Y(_03749_));
 sky130_fd_sc_hs__a21boi_1 _09423_ (.A1(_03749_),
    .A2(_03748_),
    .B1_N(net3784),
    .Y(_00457_));
 sky130_fd_sc_hs__nand2_1 _09424_ (.A(net3673),
    .B(net3745),
    .Y(_03750_));
 sky130_fd_sc_hs__a21oi_1 _09425_ (.A1(net1873),
    .A2(_03750_),
    .B1(net3783),
    .Y(_00458_));
 sky130_fd_sc_hs__nand2_1 _09426_ (.A(_00221_),
    .B(\u_window_buffer.current_state[2] ),
    .Y(_03751_));
 sky130_fd_sc_hs__nor3_1 _09427_ (.A(\u_window_buffer.current_state[3] ),
    .B(_00664_),
    .C(_02177_),
    .Y(_03752_));
 sky130_fd_sc_hs__nor2_1 _09428_ (.A(\u_window_buffer.current_state[0] ),
    .B(_02178_),
    .Y(_03753_));
 sky130_fd_sc_hs__nor2_1 _09429_ (.A(_00664_),
    .B(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hs__inv_2 _09430_ (.A(net3331),
    .Y(_03755_));
 sky130_fd_sc_hs__a221oi_1 _09431_ (.A1(_03751_),
    .A2(net3379),
    .B1(_03755_),
    .B2(_00221_),
    .C1(_05774_),
    .Y(_00459_));
 sky130_fd_sc_hs__nor3_1 _09432_ (.A(_00634_),
    .B(_00651_),
    .C(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hs__a21oi_1 _09433_ (.A1(net3331),
    .A2(_00613_),
    .B1(net3782),
    .Y(_03757_));
 sky130_fd_sc_hs__buf_1 place2117 (.A(_04602_),
    .X(net2117));
 sky130_fd_sc_hs__o21ai_1 _09435_ (.A1(\u_window_buffer.move_counter[10] ),
    .A2(_03756_),
    .B1(net3292),
    .Y(_03759_));
 sky130_fd_sc_hs__a21oi_1 _09436_ (.A1(\u_window_buffer.move_counter[10] ),
    .A2(_03756_),
    .B1(_03759_),
    .Y(_00460_));
 sky130_fd_sc_hs__nor3_1 _09437_ (.A(\u_window_buffer.move_counter[2] ),
    .B(\u_window_buffer.move_counter[0] ),
    .C(\u_window_buffer.move_counter[1] ),
    .Y(_03760_));
 sky130_fd_sc_hs__nor2_1 _09438_ (.A(\u_window_buffer.move_counter[3] ),
    .B(\u_window_buffer.move_counter[4] ),
    .Y(_03761_));
 sky130_fd_sc_hs__nand2_1 _09439_ (.A(_03760_),
    .B(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hs__nor2_1 _09440_ (.A(_03762_),
    .B(_03755_),
    .Y(_03763_));
 sky130_fd_sc_hs__nor3_1 _09441_ (.A(\u_window_buffer.move_counter[5] ),
    .B(\u_window_buffer.move_counter[8] ),
    .C(_00647_),
    .Y(_03764_));
 sky130_fd_sc_hs__and2_1 _09442_ (.A(_03763_),
    .B(_03764_),
    .X(_03765_));
 sky130_fd_sc_hs__nor2_1 _09443_ (.A(\u_window_buffer.move_counter[9] ),
    .B(\u_window_buffer.move_counter[10] ),
    .Y(_03766_));
 sky130_fd_sc_hs__and2_1 _09444_ (.A(_03765_),
    .B(_03766_),
    .X(_03767_));
 sky130_fd_sc_hs__o21ai_1 _09445_ (.A1(\u_window_buffer.move_counter[11] ),
    .A2(_03767_),
    .B1(net3292),
    .Y(_03768_));
 sky130_fd_sc_hs__a21oi_1 _09446_ (.A1(\u_window_buffer.move_counter[11] ),
    .A2(_03767_),
    .B1(_03768_),
    .Y(_00461_));
 sky130_fd_sc_hs__nand3_1 _09447_ (.A(_00635_),
    .B(_00648_),
    .C(_00642_),
    .Y(_03769_));
 sky130_fd_sc_hs__nor2_1 _09448_ (.A(_03769_),
    .B(_03755_),
    .Y(_03770_));
 sky130_fd_sc_hs__o21ai_1 _09449_ (.A1(\u_window_buffer.move_counter[12] ),
    .A2(_03770_),
    .B1(net3292),
    .Y(_03771_));
 sky130_fd_sc_hs__a21oi_1 _09450_ (.A1(\u_window_buffer.move_counter[12] ),
    .A2(_03770_),
    .B1(_03771_),
    .Y(_00462_));
 sky130_fd_sc_hs__nand3b_1 _09451_ (.A_N(_03762_),
    .B(_03764_),
    .C(_03766_),
    .Y(_03772_));
 sky130_fd_sc_hs__nor3_1 _09452_ (.A(\u_window_buffer.move_counter[11] ),
    .B(\u_window_buffer.move_counter[12] ),
    .C(_03772_),
    .Y(_03773_));
 sky130_fd_sc_hs__inv_1 _09453_ (.A(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hs__nor2_1 _09454_ (.A(_03755_),
    .B(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hs__inv_1 _09455_ (.A(_03775_),
    .Y(_03776_));
 sky130_fd_sc_hs__nand2_1 _09456_ (.A(_03776_),
    .B(\u_window_buffer.move_counter[13] ),
    .Y(_03777_));
 sky130_fd_sc_hs__inv_1 _09457_ (.A(\u_window_buffer.move_counter[13] ),
    .Y(_03778_));
 sky130_fd_sc_hs__nand2_1 _09458_ (.A(_03775_),
    .B(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hs__inv_2 _09459_ (.A(_03757_),
    .Y(_03780_));
 sky130_fd_sc_hs__buf_1 place2116 (.A(_05483_),
    .X(net2116));
 sky130_fd_sc_hs__a21oi_1 _09461_ (.A1(_03777_),
    .A2(_03779_),
    .B1(_03780_),
    .Y(_00463_));
 sky130_fd_sc_hs__a21oi_1 _09462_ (.A1(_03770_),
    .A2(_00637_),
    .B1(\u_window_buffer.move_counter[14] ),
    .Y(_03782_));
 sky130_fd_sc_hs__inv_1 _09463_ (.A(\u_window_buffer.move_counter[14] ),
    .Y(_03783_));
 sky130_fd_sc_hs__inv_1 _09464_ (.A(_00637_),
    .Y(_03784_));
 sky130_fd_sc_hs__nor4_1 _09465_ (.A(_03783_),
    .B(_03784_),
    .C(_03769_),
    .D(_03755_),
    .Y(_03785_));
 sky130_fd_sc_hs__nor3_1 _09466_ (.A(_03780_),
    .B(_03782_),
    .C(_03785_),
    .Y(_00464_));
 sky130_fd_sc_hs__inv_1 _09467_ (.A(\u_window_buffer.move_counter[15] ),
    .Y(_03786_));
 sky130_fd_sc_hs__nand3_1 _09468_ (.A(_03775_),
    .B(_03778_),
    .C(_03783_),
    .Y(_03787_));
 sky130_fd_sc_hs__o21ai_1 _09469_ (.A1(_03786_),
    .A2(_03787_),
    .B1(net3292),
    .Y(_03788_));
 sky130_fd_sc_hs__a21oi_1 _09470_ (.A1(_03786_),
    .A2(_03787_),
    .B1(_03788_),
    .Y(_00465_));
 sky130_fd_sc_hs__nor2_1 _09471_ (.A(_03755_),
    .B(_00653_),
    .Y(_03789_));
 sky130_fd_sc_hs__o21ai_1 _09472_ (.A1(\u_window_buffer.move_counter[16] ),
    .A2(_03789_),
    .B1(net3292),
    .Y(_03790_));
 sky130_fd_sc_hs__a21oi_1 _09473_ (.A1(\u_window_buffer.move_counter[16] ),
    .A2(_03789_),
    .B1(_03790_),
    .Y(_00466_));
 sky130_fd_sc_hs__nand3b_1 _09474_ (.A_N(\u_window_buffer.move_counter[16] ),
    .B(_00636_),
    .C(_03778_),
    .Y(_03791_));
 sky130_fd_sc_hs__nor2_1 _09475_ (.A(_03791_),
    .B(_03776_),
    .Y(_03792_));
 sky130_fd_sc_hs__inv_1 _09476_ (.A(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hs__or2_1 _09477_ (.A(\u_window_buffer.move_counter[17] ),
    .B(_03793_),
    .X(_03794_));
 sky130_fd_sc_hs__nand2_1 _09478_ (.A(_03793_),
    .B(\u_window_buffer.move_counter[17] ),
    .Y(_03795_));
 sky130_fd_sc_hs__a21oi_1 _09479_ (.A1(_03794_),
    .A2(_03795_),
    .B1(_03780_),
    .Y(_00467_));
 sky130_fd_sc_hs__inv_1 _09480_ (.A(\u_window_buffer.move_counter[18] ),
    .Y(_03796_));
 sky130_fd_sc_hs__nor2_1 _09481_ (.A(_00632_),
    .B(_03784_),
    .Y(_03797_));
 sky130_fd_sc_hs__nand4_1 _09482_ (.A(_03756_),
    .B(_00625_),
    .C(_00636_),
    .D(_03797_),
    .Y(_03798_));
 sky130_fd_sc_hs__o21ai_1 _09483_ (.A1(_03796_),
    .A2(_03798_),
    .B1(net3292),
    .Y(_03799_));
 sky130_fd_sc_hs__a21oi_1 _09484_ (.A1(_03796_),
    .A2(_03798_),
    .B1(_03799_),
    .Y(_00468_));
 sky130_fd_sc_hs__nor2_1 _09485_ (.A(\u_window_buffer.move_counter[17] ),
    .B(\u_window_buffer.move_counter[18] ),
    .Y(_03800_));
 sky130_fd_sc_hs__inv_2 _09486_ (.A(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hs__nor3_1 _09487_ (.A(_03791_),
    .B(_03801_),
    .C(_03774_),
    .Y(_03802_));
 sky130_fd_sc_hs__nand2_1 _09488_ (.A(_03802_),
    .B(net3331),
    .Y(_03803_));
 sky130_fd_sc_hs__or2_1 _09489_ (.A(\u_window_buffer.move_counter[19] ),
    .B(_03803_),
    .X(_03804_));
 sky130_fd_sc_hs__nand2_1 _09490_ (.A(_03803_),
    .B(\u_window_buffer.move_counter[19] ),
    .Y(_03805_));
 sky130_fd_sc_hs__a21oi_1 _09491_ (.A1(_03804_),
    .A2(_03805_),
    .B1(_03780_),
    .Y(_00469_));
 sky130_fd_sc_hs__o21a_1 _09492_ (.A1(_00613_),
    .A2(_00224_),
    .B1(net3379),
    .X(_03806_));
 sky130_fd_sc_hs__a211oi_1 _09493_ (.A1(_03755_),
    .A2(_00222_),
    .B1(_05774_),
    .C1(_03806_),
    .Y(_00470_));
 sky130_fd_sc_hs__nor2_1 _09494_ (.A(_00624_),
    .B(_03798_),
    .Y(_03807_));
 sky130_fd_sc_hs__a21oi_1 _09495_ (.A1(_03807_),
    .A2(\u_window_buffer.move_counter[20] ),
    .B1(_03780_),
    .Y(_03808_));
 sky130_fd_sc_hs__o21a_1 _09496_ (.A1(\u_window_buffer.move_counter[20] ),
    .A2(_03807_),
    .B1(_03808_),
    .X(_00471_));
 sky130_fd_sc_hs__nor2_1 _09497_ (.A(\u_window_buffer.move_counter[19] ),
    .B(\u_window_buffer.move_counter[20] ),
    .Y(_03809_));
 sky130_fd_sc_hs__inv_1 _09498_ (.A(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hs__nor2_1 _09499_ (.A(_03801_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hs__nand2_1 _09500_ (.A(_03792_),
    .B(_03811_),
    .Y(_03812_));
 sky130_fd_sc_hs__or2_1 _09501_ (.A(\u_window_buffer.move_counter[21] ),
    .B(_03812_),
    .X(_03813_));
 sky130_fd_sc_hs__nand2_1 _09502_ (.A(_03812_),
    .B(\u_window_buffer.move_counter[21] ),
    .Y(_03814_));
 sky130_fd_sc_hs__a21oi_1 _09503_ (.A1(_03813_),
    .A2(_03814_),
    .B1(_03780_),
    .Y(_00472_));
 sky130_fd_sc_hs__inv_1 _09504_ (.A(_03807_),
    .Y(_03815_));
 sky130_fd_sc_hs__nor2_1 _09505_ (.A(_00617_),
    .B(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hs__o21ai_1 _09506_ (.A1(\u_window_buffer.move_counter[22] ),
    .A2(_03816_),
    .B1(net3292),
    .Y(_03817_));
 sky130_fd_sc_hs__a21oi_1 _09507_ (.A1(\u_window_buffer.move_counter[22] ),
    .A2(_03816_),
    .B1(_03817_),
    .Y(_00473_));
 sky130_fd_sc_hs__inv_1 _09508_ (.A(\u_window_buffer.move_counter[23] ),
    .Y(_03818_));
 sky130_fd_sc_hs__nor2_1 _09509_ (.A(\u_window_buffer.move_counter[21] ),
    .B(\u_window_buffer.move_counter[22] ),
    .Y(_03819_));
 sky130_fd_sc_hs__nand4_1 _09510_ (.A(_03802_),
    .B(net3331),
    .C(_03809_),
    .D(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hs__a21oi_1 _09511_ (.A1(_03820_),
    .A2(_03818_),
    .B1(_03780_),
    .Y(_03821_));
 sky130_fd_sc_hs__o21a_1 _09512_ (.A1(_03818_),
    .A2(_03820_),
    .B1(_03821_),
    .X(_00474_));
 sky130_fd_sc_hs__nand4_1 _09513_ (.A(_03789_),
    .B(_00614_),
    .C(_00616_),
    .D(_00627_),
    .Y(_03822_));
 sky130_fd_sc_hs__o21ai_1 _09514_ (.A1(_00619_),
    .A2(_03822_),
    .B1(net3292),
    .Y(_03823_));
 sky130_fd_sc_hs__a21oi_1 _09515_ (.A1(_00619_),
    .A2(_03822_),
    .B1(_03823_),
    .Y(_00475_));
 sky130_fd_sc_hs__nor4_1 _09516_ (.A(\u_window_buffer.move_counter[21] ),
    .B(\u_window_buffer.move_counter[24] ),
    .C(_00615_),
    .D(_03812_),
    .Y(_03824_));
 sky130_fd_sc_hs__o21ai_1 _09517_ (.A1(\u_window_buffer.move_counter[25] ),
    .A2(_03824_),
    .B1(net3292),
    .Y(_03825_));
 sky130_fd_sc_hs__a21oi_1 _09518_ (.A1(\u_window_buffer.move_counter[25] ),
    .A2(_03824_),
    .B1(_03825_),
    .Y(_00476_));
 sky130_fd_sc_hs__nor2_1 _09519_ (.A(\u_window_buffer.move_counter[25] ),
    .B(\u_window_buffer.move_counter[24] ),
    .Y(_03826_));
 sky130_fd_sc_hs__nand3_1 _09520_ (.A(_03816_),
    .B(_00614_),
    .C(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hs__clkinv_1 _09521_ (.A(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hs__o21ai_1 _09522_ (.A1(\u_window_buffer.move_counter[26] ),
    .A2(_03828_),
    .B1(net3292),
    .Y(_03829_));
 sky130_fd_sc_hs__a21oi_1 _09523_ (.A1(\u_window_buffer.move_counter[26] ),
    .A2(_03828_),
    .B1(_03829_),
    .Y(_00477_));
 sky130_fd_sc_hs__nand2_1 _09524_ (.A(_03824_),
    .B(_00618_),
    .Y(_03830_));
 sky130_fd_sc_hs__o21ai_1 _09525_ (.A1(_00620_),
    .A2(_03830_),
    .B1(net3292),
    .Y(_03831_));
 sky130_fd_sc_hs__a21oi_1 _09526_ (.A1(_00620_),
    .A2(_03830_),
    .B1(_03831_),
    .Y(_00478_));
 sky130_fd_sc_hs__and3_1 _09527_ (.A(_03807_),
    .B(\u_window_buffer.move_counter[28] ),
    .C(_00622_),
    .X(_03832_));
 sky130_fd_sc_hs__a21oi_1 _09528_ (.A1(_03807_),
    .A2(_00622_),
    .B1(\u_window_buffer.move_counter[28] ),
    .Y(_03833_));
 sky130_fd_sc_hs__nor3_1 _09529_ (.A(_03780_),
    .B(_03832_),
    .C(_03833_),
    .Y(_00479_));
 sky130_fd_sc_hs__nor2_1 _09530_ (.A(\u_window_buffer.move_counter[27] ),
    .B(\u_window_buffer.move_counter[28] ),
    .Y(_03834_));
 sky130_fd_sc_hs__inv_2 _09531_ (.A(_03834_),
    .Y(_03835_));
 sky130_fd_sc_hs__nor2_1 _09532_ (.A(_03835_),
    .B(_03830_),
    .Y(_03836_));
 sky130_fd_sc_hs__o21ai_1 _09533_ (.A1(\u_window_buffer.move_counter[29] ),
    .A2(_03836_),
    .B1(net3292),
    .Y(_03837_));
 sky130_fd_sc_hs__a21oi_1 _09534_ (.A1(\u_window_buffer.move_counter[29] ),
    .A2(_03836_),
    .B1(_03837_),
    .Y(_00480_));
 sky130_fd_sc_hs__nand2_1 _09535_ (.A(\u_window_buffer.move_counter[2] ),
    .B(_00223_),
    .Y(_03838_));
 sky130_fd_sc_hs__nand2_1 _09536_ (.A(_03838_),
    .B(\u_window_buffer.current_state[2] ),
    .Y(_03839_));
 sky130_fd_sc_hs__nand2_1 _09537_ (.A(net3379),
    .B(_00639_),
    .Y(_03840_));
 sky130_fd_sc_hs__a21oi_1 _09538_ (.A1(net3331),
    .A2(_03840_),
    .B1(\u_window_buffer.move_counter[2] ),
    .Y(_03841_));
 sky130_fd_sc_hs__a211oi_1 _09539_ (.A1(net3379),
    .A2(_03839_),
    .B1(_05774_),
    .C1(_03841_),
    .Y(_00481_));
 sky130_fd_sc_hs__nor3_1 _09540_ (.A(\u_window_buffer.move_counter[26] ),
    .B(\u_window_buffer.move_counter[29] ),
    .C(_03835_),
    .Y(_03842_));
 sky130_fd_sc_hs__and3_1 _09541_ (.A(_03828_),
    .B(\u_window_buffer.move_counter[30] ),
    .C(_03842_),
    .X(_03843_));
 sky130_fd_sc_hs__a21oi_1 _09542_ (.A1(_03828_),
    .A2(_03842_),
    .B1(\u_window_buffer.move_counter[30] ),
    .Y(_03844_));
 sky130_fd_sc_hs__nor3_1 _09543_ (.A(_03780_),
    .B(_03843_),
    .C(_03844_),
    .Y(_00482_));
 sky130_fd_sc_hs__a21oi_1 _09544_ (.A1(_03836_),
    .A2(_00628_),
    .B1(\u_window_buffer.move_counter[31] ),
    .Y(_03845_));
 sky130_fd_sc_hs__a31o_1 _09545_ (.A1(_03836_),
    .A2(\u_window_buffer.move_counter[31] ),
    .A3(_00628_),
    .B1(_03780_),
    .X(_03846_));
 sky130_fd_sc_hs__nor2_1 _09546_ (.A(_03845_),
    .B(_03846_),
    .Y(_00483_));
 sky130_fd_sc_hs__buf_1 place2115 (.A(_05488_),
    .X(net2115));
 sky130_fd_sc_hs__xnor2_1 _09548_ (.A(\u_window_buffer.move_counter[3] ),
    .B(_03760_),
    .Y(_03848_));
 sky130_fd_sc_hs__or2_1 _09549_ (.A(_00613_),
    .B(_03848_),
    .X(_03849_));
 sky130_fd_sc_hs__o21ai_1 _09550_ (.A1(\u_window_buffer.move_counter[3] ),
    .A2(net3331),
    .B1(net3784),
    .Y(_03850_));
 sky130_fd_sc_hs__a21oi_1 _09551_ (.A1(net3379),
    .A2(_03849_),
    .B1(_03850_),
    .Y(_00484_));
 sky130_fd_sc_hs__nor2_1 _09552_ (.A(\u_window_buffer.current_state[3] ),
    .B(_03755_),
    .Y(_03851_));
 sky130_fd_sc_hs__a21oi_1 _09553_ (.A1(_00642_),
    .A2(\u_window_buffer.move_counter[4] ),
    .B1(_00613_),
    .Y(_03852_));
 sky130_fd_sc_hs__o21ai_1 _09554_ (.A1(\u_window_buffer.move_counter[4] ),
    .A2(_00642_),
    .B1(_03852_),
    .Y(_03853_));
 sky130_fd_sc_hs__o21ai_1 _09555_ (.A1(\u_window_buffer.move_counter[4] ),
    .A2(net3331),
    .B1(net3784),
    .Y(_03854_));
 sky130_fd_sc_hs__a21oi_1 _09556_ (.A1(_03851_),
    .A2(_03853_),
    .B1(_03854_),
    .Y(_00485_));
 sky130_fd_sc_hs__o21ai_1 _09557_ (.A1(\u_window_buffer.move_counter[5] ),
    .A2(_03763_),
    .B1(net3292),
    .Y(_03855_));
 sky130_fd_sc_hs__a21oi_1 _09558_ (.A1(\u_window_buffer.move_counter[5] ),
    .A2(_03763_),
    .B1(_03855_),
    .Y(_00486_));
 sky130_fd_sc_hs__nand3_1 _09559_ (.A(net3331),
    .B(_00644_),
    .C(_00642_),
    .Y(_03856_));
 sky130_fd_sc_hs__xor2_1 _09560_ (.A(\u_window_buffer.move_counter[6] ),
    .B(_03856_),
    .X(_03857_));
 sky130_fd_sc_hs__nor2_1 _09561_ (.A(_03780_),
    .B(_03857_),
    .Y(_00487_));
 sky130_fd_sc_hs__nor3_1 _09562_ (.A(\u_window_buffer.move_counter[5] ),
    .B(\u_window_buffer.move_counter[6] ),
    .C(_03762_),
    .Y(_03858_));
 sky130_fd_sc_hs__a21oi_1 _09563_ (.A1(_03858_),
    .A2(\u_window_buffer.move_counter[7] ),
    .B1(_00613_),
    .Y(_03859_));
 sky130_fd_sc_hs__o21ai_1 _09564_ (.A1(\u_window_buffer.move_counter[7] ),
    .A2(_03858_),
    .B1(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hs__buf_1 place2114 (.A(_01742_),
    .X(net2114));
 sky130_fd_sc_hs__o21ai_1 _09566_ (.A1(\u_window_buffer.move_counter[7] ),
    .A2(net3331),
    .B1(net3784),
    .Y(_03862_));
 sky130_fd_sc_hs__a21oi_1 _09567_ (.A1(_03860_),
    .A2(net3379),
    .B1(_03862_),
    .Y(_00488_));
 sky130_fd_sc_hs__xnor2_1 _09568_ (.A(\u_window_buffer.move_counter[8] ),
    .B(_00650_),
    .Y(_03863_));
 sky130_fd_sc_hs__o21ai_1 _09569_ (.A1(_00613_),
    .A2(_03863_),
    .B1(_02178_),
    .Y(_03864_));
 sky130_fd_sc_hs__nand2_1 _09570_ (.A(_03864_),
    .B(net3331),
    .Y(_03865_));
 sky130_fd_sc_hs__nand2_1 _09571_ (.A(_03755_),
    .B(\u_window_buffer.move_counter[8] ),
    .Y(_03866_));
 sky130_fd_sc_hs__a21oi_1 _09572_ (.A1(_03865_),
    .A2(_03866_),
    .B1(net3782),
    .Y(_00489_));
 sky130_fd_sc_hs__o21ai_1 _09573_ (.A1(\u_window_buffer.move_counter[9] ),
    .A2(_03765_),
    .B1(net3292),
    .Y(_03867_));
 sky130_fd_sc_hs__a21oi_1 _09574_ (.A1(\u_window_buffer.move_counter[9] ),
    .A2(_03765_),
    .B1(_03867_),
    .Y(_00490_));
 sky130_fd_sc_hs__nand3_4 _09575_ (.A(net1848),
    .B(\u_window_buffer.next_state_is_valid_to_read ),
    .C(\u_hamming_window.rd_en_o ),
    .Y(_03868_));
 sky130_fd_sc_hs__buf_1 place2112 (.A(_01745_),
    .X(net2112));
 sky130_fd_sc_hs__buf_2 place2111 (.A(_03517_),
    .X(net2111));
 sky130_fd_sc_hs__o21ai_4 _09578_ (.A1(net3671),
    .A2(net1846),
    .B1(net3784),
    .Y(_03871_));
 sky130_fd_sc_hs__a21oi_1 _09579_ (.A1(net3671),
    .A2(net1846),
    .B1(_03871_),
    .Y(_00491_));
 sky130_fd_sc_hs__clkinv_1 _09580_ (.A(net3743),
    .Y(_03872_));
 sky130_fd_sc_hs__bufbuf_8 place2110 (.A(_04601_),
    .X(net2110));
 sky130_fd_sc_hs__clkinv_1 _09582_ (.A(net3723),
    .Y(_03874_));
 sky130_fd_sc_hs__inv_4 _09583_ (.A(\u_window_buffer.read_ptr[1] ),
    .Y(_03875_));
 sky130_fd_sc_hs__nor2_4 _09584_ (.A(_03874_),
    .B(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hs__nand2_2 _09585_ (.A(_03876_),
    .B(net3744),
    .Y(_03877_));
 sky130_fd_sc_hs__xnor2_1 _09586_ (.A(net3720),
    .B(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hs__nor2_1 _09587_ (.A(_00227_),
    .B(_00150_),
    .Y(_03879_));
 sky130_fd_sc_hs__inv_2 _09588_ (.A(_03879_),
    .Y(_03880_));
 sky130_fd_sc_hs__nor2_1 _09589_ (.A(net3723),
    .B(net3500),
    .Y(_03881_));
 sky130_fd_sc_hs__nand2_2 _09590_ (.A(net3723),
    .B(_00226_),
    .Y(_03882_));
 sky130_fd_sc_hs__inv_2 _09591_ (.A(net3441),
    .Y(_03883_));
 sky130_fd_sc_hs__nor2_1 _09592_ (.A(_03881_),
    .B(_03883_),
    .Y(_03884_));
 sky130_fd_sc_hs__nor2_2 _09593_ (.A(_03880_),
    .B(_03884_),
    .Y(_03885_));
 sky130_fd_sc_hs__inv_1 _09594_ (.A(net3722),
    .Y(_03886_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09595_ (.A(net3724),
    .Y(_03887_));
 sky130_fd_sc_hs__clkinv_2 _09596_ (.A(net3725),
    .Y(_03888_));
 sky130_fd_sc_hs__inv_1 _09597_ (.A(net3726),
    .Y(_03889_));
 sky130_fd_sc_hs__nor4_1 _09598_ (.A(_03886_),
    .B(_03887_),
    .C(_03888_),
    .D(_03889_),
    .Y(_03890_));
 sky130_fd_sc_hs__inv_1 _09599_ (.A(net3727),
    .Y(_03891_));
 sky130_fd_sc_hs__clkinv_1 _09600_ (.A(net3728),
    .Y(_03892_));
 sky130_fd_sc_hs__inv_1 _09601_ (.A(net3729),
    .Y(_03893_));
 sky130_fd_sc_hs__inv_2 _09602_ (.A(net3730),
    .Y(_03894_));
 sky130_fd_sc_hs__nor4_1 _09603_ (.A(_03891_),
    .B(_03892_),
    .C(_03893_),
    .D(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hs__nand2_1 _09604_ (.A(_03890_),
    .B(net3440),
    .Y(_03896_));
 sky130_fd_sc_hs__inv_4 _09605_ (.A(net3735),
    .Y(_03897_));
 sky130_fd_sc_hs__inv_2 _09606_ (.A(net3736),
    .Y(_03898_));
 sky130_fd_sc_hs__nor2_1 _09607_ (.A(_03897_),
    .B(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hs__nand3_1 _09608_ (.A(_03899_),
    .B(net3737),
    .C(net3738),
    .Y(_03900_));
 sky130_fd_sc_hs__inv_1 _09609_ (.A(net3717),
    .Y(_03901_));
 sky130_fd_sc_hs__inv_1 _09610_ (.A(net3718),
    .Y(_03902_));
 sky130_fd_sc_hs__nor2_4 _09611_ (.A(_03901_),
    .B(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hs__nand3_1 _09612_ (.A(_03903_),
    .B(net3719),
    .C(net3720),
    .Y(_03904_));
 sky130_fd_sc_hs__nor2_4 _09613_ (.A(_03904_),
    .B(_03877_),
    .Y(_03905_));
 sky130_fd_sc_hs__nand4_1 _09614_ (.A(net3739),
    .B(net3740),
    .C(net3741),
    .D(net3742),
    .Y(_03906_));
 sky130_fd_sc_hs__inv_1 _09615_ (.A(net3714),
    .Y(_03907_));
 sky130_fd_sc_hs__nor2_1 _09616_ (.A(_03872_),
    .B(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hs__and2_1 _09617_ (.A(net3715),
    .B(net3716),
    .X(_03909_));
 sky130_fd_sc_hs__nand2_1 _09618_ (.A(_03908_),
    .B(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hs__nor2_1 _09619_ (.A(_03906_),
    .B(_03910_),
    .Y(_03911_));
 sky130_fd_sc_hs__nand2_1 _09620_ (.A(_03905_),
    .B(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hs__nor2_2 _09621_ (.A(_03900_),
    .B(net3289),
    .Y(_03913_));
 sky130_fd_sc_hs__inv_1 _09622_ (.A(net3733),
    .Y(_03914_));
 sky130_fd_sc_hs__inv_4 _09623_ (.A(net3734),
    .Y(_03915_));
 sky130_fd_sc_hs__nor2_1 _09624_ (.A(_03914_),
    .B(_03915_),
    .Y(_03916_));
 sky130_fd_sc_hs__inv_1 _09625_ (.A(net3731),
    .Y(_03917_));
 sky130_fd_sc_hs__inv_1 _09626_ (.A(net3732),
    .Y(_03918_));
 sky130_fd_sc_hs__nor2_1 _09627_ (.A(_03917_),
    .B(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hs__nand3_1 _09628_ (.A(_03913_),
    .B(net3436),
    .C(_03919_),
    .Y(_03920_));
 sky130_fd_sc_hs__nor2_1 _09629_ (.A(_03896_),
    .B(net3212),
    .Y(_03921_));
 sky130_fd_sc_hs__or2_1 _09630_ (.A(net3721),
    .B(_03921_),
    .X(_03922_));
 sky130_fd_sc_hs__nand2_1 _09631_ (.A(_03921_),
    .B(net3721),
    .Y(_03923_));
 sky130_fd_sc_hs__nand2_1 _09632_ (.A(_03922_),
    .B(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hs__buf_1 place2109 (.A(_04603_),
    .X(net2109));
 sky130_fd_sc_hs__nor2_1 _09634_ (.A(net3291),
    .B(net3075),
    .Y(_03926_));
 sky130_fd_sc_hs__xnor2_1 _09635_ (.A(net3330),
    .B(_03926_),
    .Y(_03927_));
 sky130_fd_sc_hs__nand2_1 _09636_ (.A(_03927_),
    .B(net3377),
    .Y(_03928_));
 sky130_fd_sc_hs__clkdlyinv3sd2_1 _09637_ (.A(net3740),
    .Y(_03929_));
 sky130_fd_sc_hs__inv_1 _09638_ (.A(net3741),
    .Y(_03930_));
 sky130_fd_sc_hs__nor2_2 _09639_ (.A(_03929_),
    .B(_03930_),
    .Y(_03931_));
 sky130_fd_sc_hs__nand3_1 _09640_ (.A(_03931_),
    .B(net3738),
    .C(net3739),
    .Y(_03932_));
 sky130_fd_sc_hs__inv_1 _09641_ (.A(net3716),
    .Y(_03933_));
 sky130_fd_sc_hs__nand2_1 _09642_ (.A(net3714),
    .B(net3715),
    .Y(_03934_));
 sky130_fd_sc_hs__nand2_1 _09643_ (.A(net3719),
    .B(net3720),
    .Y(_03935_));
 sky130_fd_sc_hs__nor3_4 _09644_ (.A(net3603),
    .B(net3602),
    .C(net3578),
    .Y(_03936_));
 sky130_fd_sc_hs__nand3_2 _09645_ (.A(_03936_),
    .B(net3744),
    .C(net3718),
    .Y(_03937_));
 sky130_fd_sc_hs__nor4_2 _09646_ (.A(_03933_),
    .B(net3590),
    .C(net3579),
    .D(_03937_),
    .Y(_03938_));
 sky130_fd_sc_hs__inv_1 _09647_ (.A(net3742),
    .Y(_03939_));
 sky130_fd_sc_hs__nor2_1 _09648_ (.A(_03939_),
    .B(net3604),
    .Y(_03940_));
 sky130_fd_sc_hs__nand2_1 _09649_ (.A(net3328),
    .B(net3433),
    .Y(_03941_));
 sky130_fd_sc_hs__nor2_1 _09650_ (.A(net3375),
    .B(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hs__nand2_1 _09651_ (.A(_03942_),
    .B(net3737),
    .Y(_03943_));
 sky130_fd_sc_hs__xnor2_1 _09652_ (.A(net3736),
    .B(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hs__inv_1 _09653_ (.A(net3165),
    .Y(_03945_));
 sky130_fd_sc_hs__nand2_1 _09654_ (.A(net3438),
    .B(net3588),
    .Y(_03946_));
 sky130_fd_sc_hs__nand3_1 _09655_ (.A(net3437),
    .B(net3741),
    .C(net3742),
    .Y(_03947_));
 sky130_fd_sc_hs__nand2_1 _09656_ (.A(_03936_),
    .B(net3744),
    .Y(_03948_));
 sky130_fd_sc_hs__nor3_2 _09657_ (.A(_03946_),
    .B(_03947_),
    .C(net3374),
    .Y(_03949_));
 sky130_fd_sc_hs__xnor2_2 _09658_ (.A(net3740),
    .B(_03949_),
    .Y(_03950_));
 sky130_fd_sc_hs__inv_1 _09659_ (.A(net3739),
    .Y(_03951_));
 sky130_fd_sc_hs__nor2_4 _09660_ (.A(_03935_),
    .B(_03882_),
    .Y(_03952_));
 sky130_fd_sc_hs__nand3_2 _09661_ (.A(_03952_),
    .B(_03903_),
    .C(net3716),
    .Y(_03953_));
 sky130_fd_sc_hs__nor2_2 _09662_ (.A(_03934_),
    .B(_03953_),
    .Y(_03954_));
 sky130_fd_sc_hs__nand3_1 _09663_ (.A(net3287),
    .B(net3433),
    .C(net3434),
    .Y(_03955_));
 sky130_fd_sc_hs__xnor2_1 _09664_ (.A(_03951_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hs__nand2_1 _09665_ (.A(_03950_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hs__nand2_1 _09666_ (.A(_03954_),
    .B(_03940_),
    .Y(_03958_));
 sky130_fd_sc_hs__xnor2_1 _09667_ (.A(net3741),
    .B(net3255),
    .Y(_03959_));
 sky130_fd_sc_hs__nand2_1 _09668_ (.A(net3328),
    .B(net3743),
    .Y(_03960_));
 sky130_fd_sc_hs__a22oi_1 _09669_ (.A1(net3433),
    .A2(net3328),
    .B1(_03960_),
    .B2(net3577),
    .Y(_03961_));
 sky130_fd_sc_hs__nor2_1 _09670_ (.A(_03959_),
    .B(_03961_),
    .Y(_03962_));
 sky130_fd_sc_hs__xnor2_1 _09671_ (.A(net3718),
    .B(_03948_),
    .Y(_03963_));
 sky130_fd_sc_hs__a21oi_1 _09672_ (.A1(net3376),
    .A2(net3720),
    .B1(net3719),
    .Y(_03964_));
 sky130_fd_sc_hs__nor2_1 _09673_ (.A(net3373),
    .B(_03964_),
    .Y(_03965_));
 sky130_fd_sc_hs__nor3b_1 _09674_ (.A(_03965_),
    .B(_03878_),
    .C_N(_03885_),
    .Y(_03966_));
 sky130_fd_sc_hs__nand2_1 _09675_ (.A(net3373),
    .B(net3718),
    .Y(_03967_));
 sky130_fd_sc_hs__xnor2_1 _09676_ (.A(net3590),
    .B(_03967_),
    .Y(_03968_));
 sky130_fd_sc_hs__nand2_1 _09677_ (.A(net3251),
    .B(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hs__nor2_2 _09678_ (.A(net3326),
    .B(_03969_),
    .Y(_03970_));
 sky130_fd_sc_hs__xnor2_1 _09679_ (.A(net3715),
    .B(net3327),
    .Y(_03971_));
 sky130_fd_sc_hs__nor2_1 _09680_ (.A(net3716),
    .B(_03905_),
    .Y(_03972_));
 sky130_fd_sc_hs__nor3_1 _09681_ (.A(net3580),
    .B(net3590),
    .C(_03937_),
    .Y(_03973_));
 sky130_fd_sc_hs__nor2_1 _09682_ (.A(_03972_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hs__nor2_1 _09683_ (.A(_03971_),
    .B(_03974_),
    .Y(_03975_));
 sky130_fd_sc_hs__nand2_1 _09684_ (.A(_03970_),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hs__a21oi_1 _09685_ (.A1(net3324),
    .A2(net3715),
    .B1(net3714),
    .Y(_03977_));
 sky130_fd_sc_hs__or2_1 _09686_ (.A(net3328),
    .B(_03977_),
    .X(_03978_));
 sky130_fd_sc_hs__xnor2_1 _09687_ (.A(net3743),
    .B(net3287),
    .Y(_03979_));
 sky130_fd_sc_hs__nand2_1 _09688_ (.A(_03978_),
    .B(_03979_),
    .Y(_03980_));
 sky130_fd_sc_hs__nor2_2 _09689_ (.A(_03976_),
    .B(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hs__nand2_1 _09690_ (.A(_03962_),
    .B(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hs__nor2_2 _09691_ (.A(_03957_),
    .B(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hs__inv_1 _09692_ (.A(net3738),
    .Y(_03984_));
 sky130_fd_sc_hs__xnor2_1 _09693_ (.A(_03984_),
    .B(net3290),
    .Y(_03985_));
 sky130_fd_sc_hs__inv_1 _09694_ (.A(net3249),
    .Y(_03986_));
 sky130_fd_sc_hs__nor2_2 _09695_ (.A(_03932_),
    .B(_03958_),
    .Y(_03987_));
 sky130_fd_sc_hs__nor2_1 _09696_ (.A(net3737),
    .B(net3207),
    .Y(_03988_));
 sky130_fd_sc_hs__inv_1 _09697_ (.A(net3737),
    .Y(_03989_));
 sky130_fd_sc_hs__inv_2 _09698_ (.A(net3207),
    .Y(_03990_));
 sky130_fd_sc_hs__nor2_2 _09699_ (.A(net3574),
    .B(_03990_),
    .Y(_03991_));
 sky130_fd_sc_hs__nor2_1 _09700_ (.A(_03988_),
    .B(net3119),
    .Y(_03992_));
 sky130_fd_sc_hs__nor2_1 _09701_ (.A(_03986_),
    .B(net3071),
    .Y(_03993_));
 sky130_fd_sc_hs__nand2_2 _09702_ (.A(_03983_),
    .B(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hs__inv_2 _09703_ (.A(_03924_),
    .Y(_03995_));
 sky130_fd_sc_hs__buf_1 place2106 (.A(net5087),
    .X(net2106));
 sky130_fd_sc_hs__nand2_1 _09705_ (.A(net2953),
    .B(net3023),
    .Y(_03997_));
 sky130_fd_sc_hs__xnor2_1 _09706_ (.A(net3121),
    .B(_03997_),
    .Y(_03998_));
 sky130_fd_sc_hs__inv_1 _09707_ (.A(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hs__nor2_1 _09708_ (.A(_03894_),
    .B(_03917_),
    .Y(_04000_));
 sky130_fd_sc_hs__clkinv_2 _09709_ (.A(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hs__inv_1 _09710_ (.A(_03899_),
    .Y(_04002_));
 sky130_fd_sc_hs__nor3_1 _09711_ (.A(_03915_),
    .B(_03989_),
    .C(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hs__nor2_1 _09712_ (.A(_03918_),
    .B(_03914_),
    .Y(_04004_));
 sky130_fd_sc_hs__nand3_1 _09713_ (.A(_03987_),
    .B(net3321),
    .C(_04004_),
    .Y(_04005_));
 sky130_fd_sc_hs__nor2_2 _09714_ (.A(_04001_),
    .B(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hs__nor2_1 _09715_ (.A(net3595),
    .B(net3594),
    .Y(_04007_));
 sky130_fd_sc_hs__and2_2 _09716_ (.A(_04006_),
    .B(_04007_),
    .X(_04008_));
 sky130_fd_sc_hs__nand2_1 _09717_ (.A(net3726),
    .B(net3727),
    .Y(_04009_));
 sky130_fd_sc_hs__nor3_1 _09718_ (.A(net3600),
    .B(net3598),
    .C(net3573),
    .Y(_04010_));
 sky130_fd_sc_hs__nand2_1 _09719_ (.A(net3070),
    .B(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hs__xnor2_1 _09720_ (.A(net3722),
    .B(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hs__nor3b_4 _09721_ (.A(net3289),
    .B(_03900_),
    .C_N(_03916_),
    .Y(_04013_));
 sky130_fd_sc_hs__nand4_2 _09722_ (.A(net3435),
    .B(net3729),
    .C(net3730),
    .D(_04013_),
    .Y(_04014_));
 sky130_fd_sc_hs__xnor2_2 _09723_ (.A(_04014_),
    .B(net3595),
    .Y(_04015_));
 sky130_fd_sc_hs__xnor2_1 _09724_ (.A(net3729),
    .B(_04006_),
    .Y(_04016_));
 sky130_fd_sc_hs__and2_2 _09725_ (.A(_04015_),
    .B(_04016_),
    .X(_04017_));
 sky130_fd_sc_hs__xnor2_1 _09726_ (.A(net3730),
    .B(net3212),
    .Y(_04018_));
 sky130_fd_sc_hs__xnor2_1 _09727_ (.A(net3731),
    .B(net3162),
    .Y(_04019_));
 sky130_fd_sc_hs__nor2_2 _09728_ (.A(_04018_),
    .B(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hs__nand2_1 _09729_ (.A(_04017_),
    .B(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hs__nor2b_1 _09730_ (.A(_03920_),
    .B_N(net3439),
    .Y(_04022_));
 sky130_fd_sc_hs__xnor2_1 _09731_ (.A(net3726),
    .B(_04022_),
    .Y(_04023_));
 sky130_fd_sc_hs__inv_1 _09732_ (.A(_04023_),
    .Y(_04024_));
 sky130_fd_sc_hs__xnor2_1 _09733_ (.A(net3727),
    .B(_04008_),
    .Y(_04025_));
 sky130_fd_sc_hs__inv_1 _09734_ (.A(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hs__nor2_2 _09735_ (.A(_04024_),
    .B(_04026_),
    .Y(_04027_));
 sky130_fd_sc_hs__nor2_1 _09736_ (.A(_03888_),
    .B(_04009_),
    .Y(_04028_));
 sky130_fd_sc_hs__nand3b_1 _09737_ (.A_N(_04014_),
    .B(net3728),
    .C(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hs__xnor2_1 _09738_ (.A(net3600),
    .B(_04029_),
    .Y(_04030_));
 sky130_fd_sc_hs__nand2_1 _09739_ (.A(net3323),
    .B(net3432),
    .Y(_04031_));
 sky130_fd_sc_hs__nor3_4 _09740_ (.A(net3372),
    .B(_04031_),
    .C(_03990_),
    .Y(_04032_));
 sky130_fd_sc_hs__nand3b_1 _09741_ (.A_N(_04009_),
    .B(_04032_),
    .C(net3431),
    .Y(_04033_));
 sky130_fd_sc_hs__xnor2_2 _09742_ (.A(net3598),
    .B(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hs__nand3_1 _09743_ (.A(_04027_),
    .B(net3115),
    .C(_04034_),
    .Y(_04035_));
 sky130_fd_sc_hs__nor2_2 _09744_ (.A(_04021_),
    .B(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hs__nor2_1 _09745_ (.A(net3441),
    .B(_03878_),
    .Y(_04037_));
 sky130_fd_sc_hs__inv_1 _09746_ (.A(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hs__nor3_2 _09747_ (.A(net3286),
    .B(_03963_),
    .C(_04038_),
    .Y(_04039_));
 sky130_fd_sc_hs__xnor2_1 _09748_ (.A(net3585),
    .B(net3256),
    .Y(_04040_));
 sky130_fd_sc_hs__nand2_1 _09749_ (.A(_03991_),
    .B(net3736),
    .Y(_04041_));
 sky130_fd_sc_hs__xnor2_2 _09750_ (.A(_04041_),
    .B(net3592),
    .Y(_04042_));
 sky130_fd_sc_hs__and2b_2 _09751_ (.A_N(_04040_),
    .B(_04042_),
    .X(_04043_));
 sky130_fd_sc_hs__nand2_1 _09752_ (.A(net3207),
    .B(net3322),
    .Y(_04044_));
 sky130_fd_sc_hs__xnor2_1 _09753_ (.A(net3733),
    .B(_04044_),
    .Y(_04045_));
 sky130_fd_sc_hs__inv_1 _09754_ (.A(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hs__xnor2_1 _09755_ (.A(net3732),
    .B(net3248),
    .Y(_04047_));
 sky130_fd_sc_hs__nand3_1 _09756_ (.A(_04043_),
    .B(_04046_),
    .C(_04047_),
    .Y(_04048_));
 sky130_fd_sc_hs__nor2_2 _09757_ (.A(_03992_),
    .B(_03944_),
    .Y(_04049_));
 sky130_fd_sc_hs__nand3_2 _09758_ (.A(_04049_),
    .B(net3211),
    .C(net3249),
    .Y(_04050_));
 sky130_fd_sc_hs__nor2_2 _09759_ (.A(_04048_),
    .B(_04050_),
    .Y(_04051_));
 sky130_fd_sc_hs__inv_1 _09760_ (.A(_03979_),
    .Y(_04052_));
 sky130_fd_sc_hs__or2_1 _09761_ (.A(_04052_),
    .B(net3253),
    .X(_04053_));
 sky130_fd_sc_hs__inv_1 _09762_ (.A(_03950_),
    .Y(_04054_));
 sky130_fd_sc_hs__nor2_1 _09763_ (.A(_03959_),
    .B(_04054_),
    .Y(_04055_));
 sky130_fd_sc_hs__clkinv_2 _09764_ (.A(_04055_),
    .Y(_04056_));
 sky130_fd_sc_hs__inv_1 _09765_ (.A(_03978_),
    .Y(_04057_));
 sky130_fd_sc_hs__nor2_1 _09766_ (.A(net3284),
    .B(_04057_),
    .Y(_04058_));
 sky130_fd_sc_hs__nand3b_1 _09767_ (.A_N(net3250),
    .B(_04058_),
    .C(net3285),
    .Y(_04059_));
 sky130_fd_sc_hs__nor3_2 _09768_ (.A(_04053_),
    .B(_04056_),
    .C(_04059_),
    .Y(_04060_));
 sky130_fd_sc_hs__nand4_2 _09769_ (.A(net3206),
    .B(_04036_),
    .C(_04051_),
    .D(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hs__xnor2_1 _09770_ (.A(_04012_),
    .B(_04061_),
    .Y(_04062_));
 sky130_fd_sc_hs__nand2_1 _09771_ (.A(_04062_),
    .B(_03995_),
    .Y(_04063_));
 sky130_fd_sc_hs__inv_1 _09772_ (.A(_04012_),
    .Y(_04064_));
 sky130_fd_sc_hs__nand2_1 _09773_ (.A(_04064_),
    .B(net3073),
    .Y(_04065_));
 sky130_fd_sc_hs__nand3_1 _09774_ (.A(_04064_),
    .B(net3116),
    .C(_03995_),
    .Y(_04066_));
 sky130_fd_sc_hs__nand2_1 _09775_ (.A(_03945_),
    .B(net3019),
    .Y(_04067_));
 sky130_fd_sc_hs__nor2_4 _09776_ (.A(_03994_),
    .B(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hs__inv_1 _09777_ (.A(net3118),
    .Y(_04069_));
 sky130_fd_sc_hs__nor2_1 _09778_ (.A(net3204),
    .B(_04045_),
    .Y(_04070_));
 sky130_fd_sc_hs__and3_1 _09779_ (.A(_04069_),
    .B(net3203),
    .C(_04070_),
    .X(_04071_));
 sky130_fd_sc_hs__nand2_2 _09780_ (.A(_04068_),
    .B(_04071_),
    .Y(_04072_));
 sky130_fd_sc_hs__nor2_4 _09781_ (.A(net3160),
    .B(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hs__inv_1 _09782_ (.A(net3020),
    .Y(_04074_));
 sky130_fd_sc_hs__nor2_1 _09783_ (.A(net3066),
    .B(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hs__nand4_2 _09784_ (.A(_04073_),
    .B(net3021),
    .C(net3022),
    .D(_04075_),
    .Y(_04076_));
 sky130_fd_sc_hs__nor2_2 _09785_ (.A(_04066_),
    .B(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hs__nand3_1 _09786_ (.A(_04063_),
    .B(_04065_),
    .C(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hs__nand2_1 _09787_ (.A(_04046_),
    .B(_04047_),
    .Y(_04079_));
 sky130_fd_sc_hs__nand2_1 _09788_ (.A(_04027_),
    .B(_04017_),
    .Y(_04080_));
 sky130_fd_sc_hs__nor3b_1 _09789_ (.A(_04079_),
    .B(_04080_),
    .C_N(net3068),
    .Y(_04081_));
 sky130_fd_sc_hs__inv_1 _09790_ (.A(net3205),
    .Y(_04082_));
 sky130_fd_sc_hs__nor3b_4 _09791_ (.A(net3250),
    .B(_04082_),
    .C_N(net3285),
    .Y(_04083_));
 sky130_fd_sc_hs__nand2_1 _09792_ (.A(_04083_),
    .B(net3157),
    .Y(_04084_));
 sky130_fd_sc_hs__nor2_1 _09793_ (.A(net3159),
    .B(net3063),
    .Y(_04085_));
 sky130_fd_sc_hs__nand2_1 _09794_ (.A(net3211),
    .B(net3249),
    .Y(_04086_));
 sky130_fd_sc_hs__nand2_1 _09795_ (.A(net3018),
    .B(net2978),
    .Y(_04087_));
 sky130_fd_sc_hs__nor3_2 _09796_ (.A(_04086_),
    .B(net3113),
    .C(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hs__nand3_1 _09797_ (.A(net2908),
    .B(net3016),
    .C(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hs__nand2_1 _09798_ (.A(_04089_),
    .B(net2977),
    .Y(_04090_));
 sky130_fd_sc_hs__nand4_1 _09799_ (.A(net2908),
    .B(net3016),
    .C(net3020),
    .D(_04088_),
    .Y(_04091_));
 sky130_fd_sc_hs__nand2_1 _09800_ (.A(_04090_),
    .B(_04091_),
    .Y(_04092_));
 sky130_fd_sc_hs__nand2_1 _09801_ (.A(_04092_),
    .B(_03995_),
    .Y(_04093_));
 sky130_fd_sc_hs__o21ai_1 _09802_ (.A1(_03995_),
    .A2(net2977),
    .B1(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hs__nor3_1 _09803_ (.A(net3159),
    .B(net3113),
    .C(_04050_),
    .Y(_04095_));
 sky130_fd_sc_hs__nor2_1 _09804_ (.A(net2980),
    .B(_04048_),
    .Y(_04096_));
 sky130_fd_sc_hs__nand3b_1 _09805_ (.A_N(net3063),
    .B(_04095_),
    .C(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hs__xnor2_1 _09806_ (.A(net2979),
    .B(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hs__nand2_1 _09807_ (.A(_04098_),
    .B(_03995_),
    .Y(_04099_));
 sky130_fd_sc_hs__nand2_1 _09808_ (.A(net3021),
    .B(net3073),
    .Y(_04100_));
 sky130_fd_sc_hs__nand2_1 _09809_ (.A(_04099_),
    .B(_04100_),
    .Y(_04101_));
 sky130_fd_sc_hs__nand3_1 _09810_ (.A(_04073_),
    .B(net3021),
    .C(net3022),
    .Y(_04102_));
 sky130_fd_sc_hs__nand2_1 _09811_ (.A(_04102_),
    .B(_03995_),
    .Y(_04103_));
 sky130_fd_sc_hs__xnor2_1 _09812_ (.A(net3117),
    .B(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hs__nand4_1 _09813_ (.A(_04078_),
    .B(_04094_),
    .C(_04101_),
    .D(_04104_),
    .Y(_04105_));
 sky130_fd_sc_hs__nand2_1 _09814_ (.A(_04063_),
    .B(_04065_),
    .Y(_04106_));
 sky130_fd_sc_hs__nand2_1 _09815_ (.A(_04076_),
    .B(_03995_),
    .Y(_04107_));
 sky130_fd_sc_hs__xnor2_1 _09816_ (.A(net3116),
    .B(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hs__nor2_1 _09817_ (.A(_04106_),
    .B(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hs__nand2_1 _09818_ (.A(_04109_),
    .B(_04105_),
    .Y(_04110_));
 sky130_fd_sc_hs__nand2_1 _09819_ (.A(net2845),
    .B(net2848),
    .Y(_04111_));
 sky130_fd_sc_hs__nand3_1 _09820_ (.A(net2801),
    .B(net2846),
    .C(net2826),
    .Y(_04112_));
 sky130_fd_sc_hs__or3_1 _09821_ (.A(net2845),
    .B(net2829),
    .C(net2828),
    .X(_04113_));
 sky130_fd_sc_hs__nand2_2 _09822_ (.A(_04112_),
    .B(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hs__a21oi_1 _09823_ (.A1(net2881),
    .A2(net3069),
    .B1(net3074),
    .Y(_04115_));
 sky130_fd_sc_hs__xnor2_1 _09824_ (.A(net3161),
    .B(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hs__inv_1 _09825_ (.A(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hs__nand2_1 _09826_ (.A(net2833),
    .B(net2832),
    .Y(_04118_));
 sky130_fd_sc_hs__inv_1 _09827_ (.A(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hs__nand3_2 _09828_ (.A(_04114_),
    .B(_04117_),
    .C(_04119_),
    .Y(_04120_));
 sky130_fd_sc_hs__inv_1 _09829_ (.A(net2833),
    .Y(_04121_));
 sky130_fd_sc_hs__or2_1 _09830_ (.A(net2818),
    .B(_04121_),
    .X(_04122_));
 sky130_fd_sc_hs__nand2_2 _09831_ (.A(_04110_),
    .B(_04111_),
    .Y(_04123_));
 sky130_fd_sc_hs__nor3_2 _09832_ (.A(net2828),
    .B(_04122_),
    .C(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hs__nand2_2 _09833_ (.A(_04120_),
    .B(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hs__nor3_4 _09834_ (.A(net2830),
    .B(net2848),
    .C(_04123_),
    .Y(_04126_));
 sky130_fd_sc_hs__inv_1 _09835_ (.A(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hs__nand2_1 _09836_ (.A(_04125_),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hs__nand2_2 _09837_ (.A(_04128_),
    .B(net2825),
    .Y(_04129_));
 sky130_fd_sc_hs__nand3_1 _09838_ (.A(_04125_),
    .B(net2844),
    .C(_04127_),
    .Y(_04130_));
 sky130_fd_sc_hs__nand3b_1 _09839_ (.A_N(net3210),
    .B(net3016),
    .C(net3288),
    .Y(_04131_));
 sky130_fd_sc_hs__nor3b_1 _09840_ (.A(net3155),
    .B(_04131_),
    .C_N(net3018),
    .Y(_04132_));
 sky130_fd_sc_hs__a21oi_1 _09841_ (.A1(net2951),
    .A2(net2978),
    .B1(net3074),
    .Y(_04133_));
 sky130_fd_sc_hs__a21oi_1 _09842_ (.A1(net3025),
    .A2(net3017),
    .B1(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hs__o21ai_1 _09843_ (.A1(net3074),
    .A2(net3067),
    .B1(_04134_),
    .Y(_04135_));
 sky130_fd_sc_hs__xnor2_1 _09844_ (.A(net3069),
    .B(_04135_),
    .Y(_04136_));
 sky130_fd_sc_hs__inv_1 _09845_ (.A(_04136_),
    .Y(_04137_));
 sky130_fd_sc_hs__nand4_2 _09846_ (.A(_04129_),
    .B(_04130_),
    .C(_04137_),
    .D(net2788),
    .Y(_04138_));
 sky130_fd_sc_hs__nand2_2 _09847_ (.A(_04123_),
    .B(net2846),
    .Y(_04139_));
 sky130_fd_sc_hs__o21bai_1 _09848_ (.A1(net2816),
    .A2(_04139_),
    .B1_N(_04122_),
    .Y(_04140_));
 sky130_fd_sc_hs__and2_2 _09849_ (.A(_04140_),
    .B(net2827),
    .X(_04141_));
 sky130_fd_sc_hs__o21ai_1 _09850_ (.A1(_04126_),
    .A2(_04124_),
    .B1(_04120_),
    .Y(_04142_));
 sky130_fd_sc_hs__or2_1 _09851_ (.A(_04141_),
    .B(_04142_),
    .X(_04143_));
 sky130_fd_sc_hs__nand2_1 _09852_ (.A(_04142_),
    .B(_04141_),
    .Y(_04144_));
 sky130_fd_sc_hs__nand2_1 _09853_ (.A(_04143_),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hs__xnor2_1 _09854_ (.A(_04119_),
    .B(_04139_),
    .Y(_04146_));
 sky130_fd_sc_hs__nand2_1 _09855_ (.A(net2787),
    .B(net2825),
    .Y(_04147_));
 sky130_fd_sc_hs__nand2_1 _09856_ (.A(_04146_),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hs__inv_1 _09857_ (.A(net2847),
    .Y(_04149_));
 sky130_fd_sc_hs__o21ai_1 _09858_ (.A1(net2831),
    .A2(net2828),
    .B1(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hs__nand4_1 _09859_ (.A(_04139_),
    .B(_04150_),
    .C(net2824),
    .D(net2817),
    .Y(_04151_));
 sky130_fd_sc_hs__nand2_1 _09860_ (.A(_04148_),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hs__nand2_1 _09861_ (.A(_04152_),
    .B(_04128_),
    .Y(_04153_));
 sky130_fd_sc_hs__nand3_1 _09862_ (.A(_04125_),
    .B(_04127_),
    .C(_04146_),
    .Y(_04154_));
 sky130_fd_sc_hs__nand2_1 _09863_ (.A(_04153_),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hs__nor2_4 _09864_ (.A(_04155_),
    .B(_04145_),
    .Y(_04156_));
 sky130_fd_sc_hs__nand2_2 _09865_ (.A(_04138_),
    .B(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hs__nor2_1 _09866_ (.A(net2828),
    .B(net2794),
    .Y(_04158_));
 sky130_fd_sc_hs__o21bai_1 _09867_ (.A1(net2768),
    .A2(_04142_),
    .B1_N(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hs__and2_2 _09868_ (.A(_04159_),
    .B(net2769),
    .X(_04160_));
 sky130_fd_sc_hs__inv_1 _09869_ (.A(_04160_),
    .Y(_04161_));
 sky130_fd_sc_hs__nand2_2 _09870_ (.A(_04157_),
    .B(_04161_),
    .Y(_04162_));
 sky130_fd_sc_hs__nand2_1 _09871_ (.A(_04162_),
    .B(net2843),
    .Y(_04163_));
 sky130_fd_sc_hs__nand3_1 _09872_ (.A(_04157_),
    .B(net2860),
    .C(_04161_),
    .Y(_04164_));
 sky130_fd_sc_hs__nand2_1 _09873_ (.A(net2909),
    .B(net3025),
    .Y(_04165_));
 sky130_fd_sc_hs__xnor2_1 _09874_ (.A(net3160),
    .B(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hs__inv_1 _09875_ (.A(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hs__and2_1 _09876_ (.A(_04129_),
    .B(net2758),
    .X(_04168_));
 sky130_fd_sc_hs__nand4_2 _09877_ (.A(_04163_),
    .B(_04164_),
    .C(_04167_),
    .D(net2744),
    .Y(_04169_));
 sky130_fd_sc_hs__xnor2_1 _09878_ (.A(net2788),
    .B(_04129_),
    .Y(_04170_));
 sky130_fd_sc_hs__nand2_1 _09879_ (.A(_04168_),
    .B(net2843),
    .Y(_04171_));
 sky130_fd_sc_hs__nand2_1 _09880_ (.A(_04170_),
    .B(_04171_),
    .Y(_04172_));
 sky130_fd_sc_hs__inv_1 _09881_ (.A(net2788),
    .Y(_04173_));
 sky130_fd_sc_hs__nand4_1 _09882_ (.A(net2751),
    .B(net2759),
    .C(_04173_),
    .D(net2843),
    .Y(_04174_));
 sky130_fd_sc_hs__nand2_1 _09883_ (.A(_04172_),
    .B(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hs__nand2_1 _09884_ (.A(_04162_),
    .B(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hs__nand3_1 _09885_ (.A(_04157_),
    .B(_04170_),
    .C(_04161_),
    .Y(_04177_));
 sky130_fd_sc_hs__nand2_2 _09886_ (.A(_04176_),
    .B(_04177_),
    .Y(_04178_));
 sky130_fd_sc_hs__o21ai_1 _09887_ (.A1(_04160_),
    .A2(net2737),
    .B1(net2746),
    .Y(_04179_));
 sky130_fd_sc_hs__nand2_1 _09888_ (.A(_04179_),
    .B(net2745),
    .Y(_04180_));
 sky130_fd_sc_hs__and2_1 _09889_ (.A(_04143_),
    .B(_04144_),
    .X(_04181_));
 sky130_fd_sc_hs__inv_1 _09890_ (.A(net2745),
    .Y(_04182_));
 sky130_fd_sc_hs__o211ai_1 _09891_ (.A1(_04181_),
    .A2(_04160_),
    .B1(_04182_),
    .C1(net2746),
    .Y(_04183_));
 sky130_fd_sc_hs__nand2_1 _09892_ (.A(_04180_),
    .B(_04183_),
    .Y(_04184_));
 sky130_fd_sc_hs__nor2_4 _09893_ (.A(_04178_),
    .B(_04184_),
    .Y(_04185_));
 sky130_fd_sc_hs__nand2_2 _09894_ (.A(_04169_),
    .B(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hs__nand3_1 _09895_ (.A(net2746),
    .B(_04182_),
    .C(_04160_),
    .Y(_04187_));
 sky130_fd_sc_hs__nand2_1 _09896_ (.A(_04187_),
    .B(net2750),
    .Y(_04188_));
 sky130_fd_sc_hs__nand2_1 _09897_ (.A(_04188_),
    .B(net2731),
    .Y(_04189_));
 sky130_fd_sc_hs__nand2_2 _09898_ (.A(_04186_),
    .B(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hs__nand2_2 _09899_ (.A(_04190_),
    .B(net2842),
    .Y(_04191_));
 sky130_fd_sc_hs__nand3_1 _09900_ (.A(_04186_),
    .B(net2859),
    .C(net2711),
    .Y(_04192_));
 sky130_fd_sc_hs__xnor2_1 _09901_ (.A(net3065),
    .B(net2907),
    .Y(_04193_));
 sky130_fd_sc_hs__inv_1 _09902_ (.A(_04193_),
    .Y(_04194_));
 sky130_fd_sc_hs__nand2_1 _09903_ (.A(net2714),
    .B(net2723),
    .Y(_04195_));
 sky130_fd_sc_hs__nor2_1 _09904_ (.A(_04194_),
    .B(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hs__nand3_2 _09905_ (.A(_04191_),
    .B(_04192_),
    .C(_04196_),
    .Y(_04197_));
 sky130_fd_sc_hs__inv_1 _09906_ (.A(_04189_),
    .Y(_04198_));
 sky130_fd_sc_hs__o211ai_1 _09907_ (.A1(_04198_),
    .A2(_04185_),
    .B1(net2704),
    .C1(net2705),
    .Y(_04199_));
 sky130_fd_sc_hs__o21ai_1 _09908_ (.A1(_04198_),
    .A2(_04185_),
    .B1(net2705),
    .Y(_04200_));
 sky130_fd_sc_hs__inv_1 _09909_ (.A(net2704),
    .Y(_04201_));
 sky130_fd_sc_hs__nand2_1 _09910_ (.A(_04200_),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hs__nand2_1 _09911_ (.A(_04199_),
    .B(_04202_),
    .Y(_04203_));
 sky130_fd_sc_hs__nand2_1 _09912_ (.A(net2751),
    .B(net2759),
    .Y(_04204_));
 sky130_fd_sc_hs__xnor2_1 _09913_ (.A(net2843),
    .B(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hs__nand2_1 _09914_ (.A(net2724),
    .B(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hs__o21ai_2 _09915_ (.A1(net2743),
    .A2(net2724),
    .B1(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hs__nand3_1 _09916_ (.A(_04163_),
    .B(_04164_),
    .C(_04167_),
    .Y(_04208_));
 sky130_fd_sc_hs__xnor2_1 _09917_ (.A(_04207_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hs__nand2_1 _09918_ (.A(_04190_),
    .B(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hs__nand3_1 _09919_ (.A(_04186_),
    .B(_04207_),
    .C(_04189_),
    .Y(_04211_));
 sky130_fd_sc_hs__and2_2 _09920_ (.A(_04210_),
    .B(_04211_),
    .X(_04212_));
 sky130_fd_sc_hs__nand3_2 _09921_ (.A(_04197_),
    .B(_04203_),
    .C(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hs__nand2_1 _09922_ (.A(net2705),
    .B(_04201_),
    .Y(_04214_));
 sky130_fd_sc_hs__o21ai_1 _09923_ (.A1(net2712),
    .A2(_04214_),
    .B1(net2713),
    .Y(_04215_));
 sky130_fd_sc_hs__nand2_1 _09924_ (.A(_04215_),
    .B(net2687),
    .Y(_04216_));
 sky130_fd_sc_hs__nand2_2 _09925_ (.A(_04213_),
    .B(_04216_),
    .Y(_04217_));
 sky130_fd_sc_hs__xnor2_1 _09926_ (.A(net2658),
    .B(net2659),
    .Y(_04218_));
 sky130_fd_sc_hs__nand2_1 _09927_ (.A(_04217_),
    .B(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hs__nand3b_1 _09928_ (.A_N(net2658),
    .B(net2647),
    .C(_04216_),
    .Y(_04220_));
 sky130_fd_sc_hs__nand2_1 _09929_ (.A(_04219_),
    .B(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hs__nand2_1 _09930_ (.A(net2664),
    .B(net2703),
    .Y(_04222_));
 sky130_fd_sc_hs__nand3b_1 _09931_ (.A_N(net2703),
    .B(net2672),
    .C(net2842),
    .Y(_04223_));
 sky130_fd_sc_hs__nand2_1 _09932_ (.A(_04222_),
    .B(_04223_),
    .Y(_04224_));
 sky130_fd_sc_hs__nand2_1 _09933_ (.A(net2663),
    .B(net2671),
    .Y(_04225_));
 sky130_fd_sc_hs__nor2_2 _09934_ (.A(net2858),
    .B(_04225_),
    .Y(_04226_));
 sky130_fd_sc_hs__xnor2_1 _09935_ (.A(_04224_),
    .B(_04226_),
    .Y(_04227_));
 sky130_fd_sc_hs__nand2_1 _09936_ (.A(_04227_),
    .B(_04217_),
    .Y(_04228_));
 sky130_fd_sc_hs__nand3b_1 _09937_ (.A_N(_04224_),
    .B(net2647),
    .C(_04216_),
    .Y(_04229_));
 sky130_fd_sc_hs__nand2_1 _09938_ (.A(_04228_),
    .B(_04229_),
    .Y(_04230_));
 sky130_fd_sc_hs__nor2_4 _09939_ (.A(_04221_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hs__nand2_1 _09940_ (.A(_04217_),
    .B(net2880),
    .Y(_04232_));
 sky130_fd_sc_hs__nand3_1 _09941_ (.A(net2646),
    .B(net2858),
    .C(_04216_),
    .Y(_04233_));
 sky130_fd_sc_hs__a21oi_1 _09942_ (.A1(net2937),
    .A2(net3064),
    .B1(net3074),
    .Y(_04234_));
 sky130_fd_sc_hs__xnor2_1 _09943_ (.A(net3203),
    .B(_04234_),
    .Y(_04235_));
 sky130_fd_sc_hs__inv_1 _09944_ (.A(_04235_),
    .Y(_04236_));
 sky130_fd_sc_hs__inv_1 _09945_ (.A(net2657),
    .Y(_04237_));
 sky130_fd_sc_hs__nand4_2 _09946_ (.A(_04232_),
    .B(_04233_),
    .C(_04236_),
    .D(_04237_),
    .Y(_04238_));
 sky130_fd_sc_hs__nand2_2 _09947_ (.A(_04231_),
    .B(_04238_),
    .Y(_04239_));
 sky130_fd_sc_hs__nand2_1 _09948_ (.A(net2659),
    .B(net2658),
    .Y(_04240_));
 sky130_fd_sc_hs__o21bai_1 _09949_ (.A1(_04216_),
    .A2(_04240_),
    .B1_N(net2662),
    .Y(_04241_));
 sky130_fd_sc_hs__nand2_1 _09950_ (.A(_04241_),
    .B(net2647),
    .Y(_04242_));
 sky130_fd_sc_hs__nand2_2 _09951_ (.A(_04239_),
    .B(net2627),
    .Y(_04243_));
 sky130_fd_sc_hs__nand2_1 _09952_ (.A(_04243_),
    .B(net2857),
    .Y(_04244_));
 sky130_fd_sc_hs__nand3_1 _09953_ (.A(_04239_),
    .B(net2879),
    .C(net2627),
    .Y(_04245_));
 sky130_fd_sc_hs__xnor2_1 _09954_ (.A(net3114),
    .B(net2936),
    .Y(_04246_));
 sky130_fd_sc_hs__and2_1 _09955_ (.A(net2628),
    .B(net2640),
    .X(_04247_));
 sky130_fd_sc_hs__nand4_1 _09956_ (.A(_04244_),
    .B(_04245_),
    .C(net2905),
    .D(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hs__nand2_1 _09957_ (.A(_04232_),
    .B(net2657),
    .Y(_04249_));
 sky130_fd_sc_hs__nand2_1 _09958_ (.A(_04217_),
    .B(net2645),
    .Y(_04250_));
 sky130_fd_sc_hs__nand2_1 _09959_ (.A(_04249_),
    .B(_04250_),
    .Y(_04251_));
 sky130_fd_sc_hs__nand2_1 _09960_ (.A(_04232_),
    .B(_04233_),
    .Y(_04252_));
 sky130_fd_sc_hs__nor2_1 _09961_ (.A(net2879),
    .B(_04252_),
    .Y(_04253_));
 sky130_fd_sc_hs__or2_1 _09962_ (.A(_04251_),
    .B(_04253_),
    .X(_04254_));
 sky130_fd_sc_hs__nand2_1 _09963_ (.A(_04253_),
    .B(_04251_),
    .Y(_04255_));
 sky130_fd_sc_hs__nand2_1 _09964_ (.A(_04254_),
    .B(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hs__nand2_1 _09965_ (.A(_04256_),
    .B(_04243_),
    .Y(_04257_));
 sky130_fd_sc_hs__nand3b_1 _09966_ (.A_N(net2614),
    .B(_04239_),
    .C(net2627),
    .Y(_04258_));
 sky130_fd_sc_hs__nand2_1 _09967_ (.A(_04257_),
    .B(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hs__inv_1 _09968_ (.A(_04242_),
    .Y(_04260_));
 sky130_fd_sc_hs__o21ai_1 _09969_ (.A1(_04260_),
    .A2(net2615),
    .B1(net2620),
    .Y(_04261_));
 sky130_fd_sc_hs__nand2_1 _09970_ (.A(_04261_),
    .B(net2621),
    .Y(_04262_));
 sky130_fd_sc_hs__and2_1 _09971_ (.A(net2629),
    .B(_04220_),
    .X(_04263_));
 sky130_fd_sc_hs__inv_1 _09972_ (.A(net2621),
    .Y(_04264_));
 sky130_fd_sc_hs__o211ai_1 _09973_ (.A1(_04263_),
    .A2(_04260_),
    .B1(_04264_),
    .C1(net2620),
    .Y(_04265_));
 sky130_fd_sc_hs__nand2_1 _09974_ (.A(_04262_),
    .B(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hs__nor2_2 _09975_ (.A(_04259_),
    .B(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hs__nand2_2 _09976_ (.A(_04248_),
    .B(_04267_),
    .Y(_04268_));
 sky130_fd_sc_hs__nand2_1 _09977_ (.A(_04265_),
    .B(net2622),
    .Y(_04269_));
 sky130_fd_sc_hs__and2_2 _09978_ (.A(_04269_),
    .B(net2611),
    .X(_04270_));
 sky130_fd_sc_hs__inv_1 _09979_ (.A(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hs__nand2_2 _09980_ (.A(_04268_),
    .B(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hs__nand2_2 _09981_ (.A(_04272_),
    .B(net2906),
    .Y(_04273_));
 sky130_fd_sc_hs__inv_1 _09982_ (.A(net2905),
    .Y(_04274_));
 sky130_fd_sc_hs__nand3_1 _09983_ (.A(_04268_),
    .B(net2878),
    .C(_04271_),
    .Y(_04275_));
 sky130_fd_sc_hs__nor2_1 _09984_ (.A(net3074),
    .B(net2937),
    .Y(_04276_));
 sky130_fd_sc_hs__xnor2_1 _09985_ (.A(net3204),
    .B(_04276_),
    .Y(_04277_));
 sky130_fd_sc_hs__nand2_1 _09986_ (.A(_04244_),
    .B(_04245_),
    .Y(_04278_));
 sky130_fd_sc_hs__inv_1 _09987_ (.A(net2582),
    .Y(_04279_));
 sky130_fd_sc_hs__nand4_1 _09988_ (.A(_04273_),
    .B(_04275_),
    .C(net2877),
    .D(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hs__nor2_2 _09989_ (.A(_04274_),
    .B(_04278_),
    .Y(_04281_));
 sky130_fd_sc_hs__xnor2_1 _09990_ (.A(net2857),
    .B(net2618),
    .Y(_04282_));
 sky130_fd_sc_hs__nand2_1 _09991_ (.A(net2602),
    .B(_04282_),
    .Y(_04283_));
 sky130_fd_sc_hs__nand3_1 _09992_ (.A(net2611),
    .B(_04247_),
    .C(net2627),
    .Y(_04284_));
 sky130_fd_sc_hs__nand2_1 _09993_ (.A(_04283_),
    .B(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hs__inv_1 _09994_ (.A(_04285_),
    .Y(_04286_));
 sky130_fd_sc_hs__nand2_1 _09995_ (.A(_04281_),
    .B(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hs__o21ai_1 _09996_ (.A1(_04274_),
    .A2(_04278_),
    .B1(_04285_),
    .Y(_04288_));
 sky130_fd_sc_hs__nand2_1 _09997_ (.A(_04287_),
    .B(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hs__nand2_1 _09998_ (.A(_04272_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hs__nand3_1 _09999_ (.A(_04268_),
    .B(net2583),
    .C(net2581),
    .Y(_04291_));
 sky130_fd_sc_hs__nand2_1 _10000_ (.A(_04290_),
    .B(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hs__o21ai_1 _10001_ (.A1(net2590),
    .A2(net2575),
    .B1(net2585),
    .Y(_04293_));
 sky130_fd_sc_hs__nand2_1 _10002_ (.A(_04293_),
    .B(net2584),
    .Y(_04294_));
 sky130_fd_sc_hs__a21oi_1 _10003_ (.A1(_04281_),
    .A2(net2619),
    .B1(net2584),
    .Y(_04295_));
 sky130_fd_sc_hs__nand2_1 _10004_ (.A(_04272_),
    .B(_04295_),
    .Y(_04296_));
 sky130_fd_sc_hs__nand2_2 _10005_ (.A(_04294_),
    .B(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hs__nor2_2 _10006_ (.A(_04292_),
    .B(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hs__nand2_2 _10007_ (.A(_04280_),
    .B(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hs__nand2_1 _10008_ (.A(_04296_),
    .B(net2591),
    .Y(_04300_));
 sky130_fd_sc_hs__nand2_1 _10009_ (.A(_04300_),
    .B(net2566),
    .Y(_04301_));
 sky130_fd_sc_hs__nand2_2 _10010_ (.A(_04299_),
    .B(_04301_),
    .Y(_04302_));
 sky130_fd_sc_hs__nand2_1 _10011_ (.A(_04302_),
    .B(net2877),
    .Y(_04303_));
 sky130_fd_sc_hs__inv_1 _10012_ (.A(net2877),
    .Y(_04304_));
 sky130_fd_sc_hs__nand3_1 _10013_ (.A(net2524),
    .B(_04304_),
    .C(_04301_),
    .Y(_04305_));
 sky130_fd_sc_hs__or2_1 _10014_ (.A(net3074),
    .B(net2952),
    .X(_04306_));
 sky130_fd_sc_hs__xnor2_1 _10015_ (.A(net3019),
    .B(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hs__nand2_1 _10016_ (.A(net2547),
    .B(net2558),
    .Y(_04308_));
 sky130_fd_sc_hs__inv_1 _10017_ (.A(net2537),
    .Y(_04309_));
 sky130_fd_sc_hs__nand4_1 _10018_ (.A(_04303_),
    .B(_04305_),
    .C(_04307_),
    .D(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hs__nand2_1 _10019_ (.A(_04273_),
    .B(net2582),
    .Y(_04311_));
 sky130_fd_sc_hs__nand2_1 _10020_ (.A(net2559),
    .B(net2573),
    .Y(_04312_));
 sky130_fd_sc_hs__and2_2 _10021_ (.A(_04311_),
    .B(_04312_),
    .X(_04313_));
 sky130_fd_sc_hs__nand3_1 _10022_ (.A(net2547),
    .B(net2558),
    .C(net2877),
    .Y(_04314_));
 sky130_fd_sc_hs__nand2_1 _10023_ (.A(_04313_),
    .B(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hs__nand4_1 _10024_ (.A(net2547),
    .B(net2558),
    .C(net2877),
    .D(net2582),
    .Y(_04316_));
 sky130_fd_sc_hs__nand2_1 _10025_ (.A(_04315_),
    .B(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hs__nand2_1 _10026_ (.A(_04302_),
    .B(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hs__nand3_1 _10027_ (.A(net2524),
    .B(_04313_),
    .C(_04301_),
    .Y(_04319_));
 sky130_fd_sc_hs__nand2_1 _10028_ (.A(_04318_),
    .B(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hs__nor2_2 _10029_ (.A(_04304_),
    .B(_04308_),
    .Y(_04321_));
 sky130_fd_sc_hs__nand3_1 _10030_ (.A(_04321_),
    .B(net2574),
    .C(net2539),
    .Y(_04322_));
 sky130_fd_sc_hs__inv_1 _10031_ (.A(net2539),
    .Y(_04323_));
 sky130_fd_sc_hs__nand2_1 _10032_ (.A(net2540),
    .B(_04323_),
    .Y(_04324_));
 sky130_fd_sc_hs__nand2_1 _10033_ (.A(_04322_),
    .B(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hs__nand2_1 _10034_ (.A(_04325_),
    .B(_04302_),
    .Y(_04326_));
 sky130_fd_sc_hs__nand3_1 _10035_ (.A(net2525),
    .B(net2539),
    .C(_04301_),
    .Y(_04327_));
 sky130_fd_sc_hs__nand2_2 _10036_ (.A(_04326_),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hs__nor2_1 _10037_ (.A(_04320_),
    .B(_04328_),
    .Y(_04329_));
 sky130_fd_sc_hs__nand2_1 _10038_ (.A(_04310_),
    .B(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hs__o21ai_1 _10039_ (.A1(_04301_),
    .A2(_04324_),
    .B1(net2538),
    .Y(_04331_));
 sky130_fd_sc_hs__and2_1 _10040_ (.A(_04331_),
    .B(net2525),
    .X(_04332_));
 sky130_fd_sc_hs__inv_1 _10041_ (.A(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hs__nand2_2 _10042_ (.A(_04330_),
    .B(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hs__nand2_2 _10043_ (.A(_04334_),
    .B(net2904),
    .Y(_04335_));
 sky130_fd_sc_hs__inv_1 _10044_ (.A(_04307_),
    .Y(_04336_));
 sky130_fd_sc_hs__nand3_1 _10045_ (.A(_04330_),
    .B(net2876),
    .C(_04333_),
    .Y(_04337_));
 sky130_fd_sc_hs__nand2_1 _10046_ (.A(_04303_),
    .B(_04305_),
    .Y(_04338_));
 sky130_fd_sc_hs__inv_1 _10047_ (.A(net2493),
    .Y(_04339_));
 sky130_fd_sc_hs__nand3_1 _10048_ (.A(_04335_),
    .B(_04337_),
    .C(_04339_),
    .Y(_04340_));
 sky130_fd_sc_hs__nor2_2 _10049_ (.A(_03999_),
    .B(_04340_),
    .Y(_04341_));
 sky130_fd_sc_hs__nand3_1 _10050_ (.A(_04334_),
    .B(net2904),
    .C(_04339_),
    .Y(_04342_));
 sky130_fd_sc_hs__a22oi_1 _10051_ (.A1(net2531),
    .A2(net2517),
    .B1(net2505),
    .B2(net2537),
    .Y(_04343_));
 sky130_fd_sc_hs__nand2_2 _10052_ (.A(_04342_),
    .B(_04343_),
    .Y(_04344_));
 sky130_fd_sc_hs__nand4_1 _10053_ (.A(_04334_),
    .B(net2904),
    .C(net2537),
    .D(_04339_),
    .Y(_04345_));
 sky130_fd_sc_hs__nor3_1 _10054_ (.A(_04336_),
    .B(net2537),
    .C(_04338_),
    .Y(_04346_));
 sky130_fd_sc_hs__nor2_1 _10055_ (.A(net2496),
    .B(_04346_),
    .Y(_04347_));
 sky130_fd_sc_hs__nand2_1 _10056_ (.A(_04334_),
    .B(_04347_),
    .Y(_04348_));
 sky130_fd_sc_hs__o21ai_1 _10057_ (.A1(_04333_),
    .A2(_04346_),
    .B1(net2496),
    .Y(_04349_));
 sky130_fd_sc_hs__and2_2 _10058_ (.A(_04348_),
    .B(_04349_),
    .X(_04350_));
 sky130_fd_sc_hs__nand3_2 _10059_ (.A(_04344_),
    .B(net2460),
    .C(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hs__nand2_1 _10060_ (.A(_04348_),
    .B(net2495),
    .Y(_04352_));
 sky130_fd_sc_hs__nand2_4 _10061_ (.A(_04352_),
    .B(net2484),
    .Y(_04353_));
 sky130_fd_sc_hs__o21ai_4 _10062_ (.A1(_04341_),
    .A2(_04351_),
    .B1(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hs__nand2_1 _10063_ (.A(_04354_),
    .B(_03999_),
    .Y(_04355_));
 sky130_fd_sc_hs__and2_1 _10064_ (.A(_04344_),
    .B(_04345_),
    .X(_04356_));
 sky130_fd_sc_hs__nand4_1 _10065_ (.A(net2462),
    .B(net2473),
    .C(_03998_),
    .D(net2489),
    .Y(_04357_));
 sky130_fd_sc_hs__nand3_2 _10066_ (.A(_04356_),
    .B(net2452),
    .C(_04357_),
    .Y(_04358_));
 sky130_fd_sc_hs__nand3_1 _10067_ (.A(_04358_),
    .B(_03998_),
    .C(_04353_),
    .Y(_04359_));
 sky130_fd_sc_hs__nand2_2 _10068_ (.A(_04355_),
    .B(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hs__inv_1 _10069_ (.A(net3072),
    .Y(_04361_));
 sky130_fd_sc_hs__o21ai_1 _10070_ (.A1(net3155),
    .A2(net2976),
    .B1(net3023),
    .Y(_04362_));
 sky130_fd_sc_hs__xnor2_1 _10071_ (.A(_04361_),
    .B(_04362_),
    .Y(_04363_));
 sky130_fd_sc_hs__nand2_1 _10072_ (.A(net2462),
    .B(net2473),
    .Y(_04364_));
 sky130_fd_sc_hs__inv_1 _10073_ (.A(net2450),
    .Y(_04365_));
 sky130_fd_sc_hs__nand3_2 _10074_ (.A(_04360_),
    .B(_04363_),
    .C(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hs__nand2_1 _10075_ (.A(_04335_),
    .B(net2494),
    .Y(_04367_));
 sky130_fd_sc_hs__nand2_1 _10076_ (.A(_04367_),
    .B(net2461),
    .Y(_04368_));
 sky130_fd_sc_hs__nor2_1 _10077_ (.A(_03999_),
    .B(_04364_),
    .Y(_04369_));
 sky130_fd_sc_hs__xnor2_1 _10078_ (.A(_04368_),
    .B(_04369_),
    .Y(_04370_));
 sky130_fd_sc_hs__nand2_1 _10079_ (.A(_04354_),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hs__inv_1 _10080_ (.A(_04368_),
    .Y(_04372_));
 sky130_fd_sc_hs__nand3_1 _10081_ (.A(_04358_),
    .B(_04353_),
    .C(_04372_),
    .Y(_04373_));
 sky130_fd_sc_hs__nand2_1 _10082_ (.A(_04371_),
    .B(_04373_),
    .Y(_04374_));
 sky130_fd_sc_hs__nand2_1 _10083_ (.A(_04344_),
    .B(_04345_),
    .Y(_04375_));
 sky130_fd_sc_hs__xnor2_1 _10084_ (.A(_04375_),
    .B(_04341_),
    .Y(_04376_));
 sky130_fd_sc_hs__nand2_1 _10085_ (.A(_04354_),
    .B(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hs__nand3_1 _10086_ (.A(_04358_),
    .B(net2443),
    .C(net2442),
    .Y(_04378_));
 sky130_fd_sc_hs__nand2_1 _10087_ (.A(_04377_),
    .B(_04378_),
    .Y(_04379_));
 sky130_fd_sc_hs__nor2_4 _10088_ (.A(_04374_),
    .B(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hs__nand2_2 _10089_ (.A(_04380_),
    .B(_04366_),
    .Y(_04381_));
 sky130_fd_sc_hs__nor2_1 _10090_ (.A(_04341_),
    .B(net2444),
    .Y(_04382_));
 sky130_fd_sc_hs__nor2_1 _10091_ (.A(_04375_),
    .B(net2445),
    .Y(_04383_));
 sky130_fd_sc_hs__inv_1 _10092_ (.A(_04353_),
    .Y(_04384_));
 sky130_fd_sc_hs__a21oi_1 _10093_ (.A1(_04383_),
    .A2(_04384_),
    .B1(net2451),
    .Y(_04385_));
 sky130_fd_sc_hs__nor2_2 _10094_ (.A(_04382_),
    .B(_04385_),
    .Y(_04386_));
 sky130_fd_sc_hs__inv_1 _10095_ (.A(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hs__nand3_1 _10096_ (.A(_04381_),
    .B(_04363_),
    .C(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hs__inv_1 _10097_ (.A(_04363_),
    .Y(_04389_));
 sky130_fd_sc_hs__o21ai_1 _10098_ (.A1(net2411),
    .A2(_04380_),
    .B1(_04389_),
    .Y(_04390_));
 sky130_fd_sc_hs__nand2_2 _10099_ (.A(_04388_),
    .B(_04390_),
    .Y(_04391_));
 sky130_fd_sc_hs__o21ai_1 _10100_ (.A1(net3164),
    .A2(net3026),
    .B1(net3023),
    .Y(_04392_));
 sky130_fd_sc_hs__xnor2_1 _10101_ (.A(net3208),
    .B(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hs__inv_1 _10102_ (.A(_04393_),
    .Y(_04394_));
 sky130_fd_sc_hs__nand3_2 _10103_ (.A(_04391_),
    .B(_04394_),
    .C(net2414),
    .Y(_04395_));
 sky130_fd_sc_hs__o21ai_1 _10104_ (.A1(_04386_),
    .A2(_04380_),
    .B1(_04366_),
    .Y(_04396_));
 sky130_fd_sc_hs__nand2_1 _10105_ (.A(_04396_),
    .B(net2413),
    .Y(_04397_));
 sky130_fd_sc_hs__and2_1 _10106_ (.A(_04377_),
    .B(_04378_),
    .X(_04398_));
 sky130_fd_sc_hs__inv_1 _10107_ (.A(net2413),
    .Y(_04399_));
 sky130_fd_sc_hs__o211ai_1 _10108_ (.A1(_04386_),
    .A2(_04398_),
    .B1(_04399_),
    .C1(_04366_),
    .Y(_04400_));
 sky130_fd_sc_hs__nand2_1 _10109_ (.A(_04397_),
    .B(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hs__nand2_1 _10110_ (.A(_04381_),
    .B(_04387_),
    .Y(_04402_));
 sky130_fd_sc_hs__xnor2_1 _10111_ (.A(_03998_),
    .B(net2450),
    .Y(_04403_));
 sky130_fd_sc_hs__nand2_1 _10112_ (.A(net2434),
    .B(_04403_),
    .Y(_04404_));
 sky130_fd_sc_hs__o21ai_1 _10113_ (.A1(net2450),
    .A2(net2434),
    .B1(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hs__nand2_1 _10114_ (.A(_04360_),
    .B(_04363_),
    .Y(_04406_));
 sky130_fd_sc_hs__xnor2_1 _10115_ (.A(_04405_),
    .B(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hs__nand2_1 _10116_ (.A(_04402_),
    .B(_04407_),
    .Y(_04408_));
 sky130_fd_sc_hs__nand3_1 _10117_ (.A(_04381_),
    .B(_04387_),
    .C(_04405_),
    .Y(_04409_));
 sky130_fd_sc_hs__nand2_2 _10118_ (.A(_04408_),
    .B(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hs__nor2_2 _10119_ (.A(_04401_),
    .B(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hs__nand2_2 _10120_ (.A(_04395_),
    .B(_04411_),
    .Y(_04412_));
 sky130_fd_sc_hs__nand2_1 _10121_ (.A(_04400_),
    .B(net2412),
    .Y(_04413_));
 sky130_fd_sc_hs__and2_1 _10122_ (.A(_04413_),
    .B(net2391),
    .X(_04414_));
 sky130_fd_sc_hs__inv_1 _10123_ (.A(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hs__nand2_2 _10124_ (.A(_04412_),
    .B(_04415_),
    .Y(_04416_));
 sky130_fd_sc_hs__nand2_2 _10125_ (.A(_04416_),
    .B(_04394_),
    .Y(_04417_));
 sky130_fd_sc_hs__nand3_1 _10126_ (.A(_04412_),
    .B(_04393_),
    .C(_04415_),
    .Y(_04418_));
 sky130_fd_sc_hs__nand2_1 _10127_ (.A(net2976),
    .B(net3023),
    .Y(_04419_));
 sky130_fd_sc_hs__xnor2_1 _10128_ (.A(net3211),
    .B(_04419_),
    .Y(_04420_));
 sky130_fd_sc_hs__nand4_2 _10129_ (.A(_04417_),
    .B(_04418_),
    .C(_04420_),
    .D(net2377),
    .Y(_04421_));
 sky130_fd_sc_hs__xnor2_1 _10130_ (.A(_04389_),
    .B(net2414),
    .Y(_04422_));
 sky130_fd_sc_hs__nand2_1 _10131_ (.A(net2385),
    .B(_04422_),
    .Y(_04423_));
 sky130_fd_sc_hs__nand3_1 _10132_ (.A(net2392),
    .B(net2400),
    .C(net2414),
    .Y(_04424_));
 sky130_fd_sc_hs__nand2_1 _10133_ (.A(_04423_),
    .B(_04424_),
    .Y(_04425_));
 sky130_fd_sc_hs__nand2_1 _10134_ (.A(net2376),
    .B(_04394_),
    .Y(_04426_));
 sky130_fd_sc_hs__xnor2_1 _10135_ (.A(_04425_),
    .B(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hs__nand2_1 _10136_ (.A(_04416_),
    .B(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hs__nand3_1 _10137_ (.A(net2350),
    .B(_04415_),
    .C(net2360),
    .Y(_04429_));
 sky130_fd_sc_hs__nand2_2 _10138_ (.A(_04428_),
    .B(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hs__o21ai_1 _10139_ (.A1(net2374),
    .A2(net2354),
    .B1(net2362),
    .Y(_04431_));
 sky130_fd_sc_hs__nand2_1 _10140_ (.A(_04431_),
    .B(net2361),
    .Y(_04432_));
 sky130_fd_sc_hs__inv_1 _10141_ (.A(net2361),
    .Y(_04433_));
 sky130_fd_sc_hs__and2_1 _10142_ (.A(net2362),
    .B(_04433_),
    .X(_04434_));
 sky130_fd_sc_hs__nand2_1 _10143_ (.A(_04416_),
    .B(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hs__nand2_2 _10144_ (.A(_04432_),
    .B(_04435_),
    .Y(_04436_));
 sky130_fd_sc_hs__nor2_4 _10145_ (.A(_04430_),
    .B(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hs__nand2_2 _10146_ (.A(_04437_),
    .B(_04421_),
    .Y(_04438_));
 sky130_fd_sc_hs__nand2_1 _10147_ (.A(net2362),
    .B(_04433_),
    .Y(_04439_));
 sky130_fd_sc_hs__o21ai_1 _10148_ (.A1(_04415_),
    .A2(_04439_),
    .B1(net2375),
    .Y(_04440_));
 sky130_fd_sc_hs__nand2_1 _10149_ (.A(_04440_),
    .B(net2349),
    .Y(_04441_));
 sky130_fd_sc_hs__nand2_2 _10150_ (.A(_04438_),
    .B(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hs__inv_1 _10151_ (.A(net2377),
    .Y(_04443_));
 sky130_fd_sc_hs__xnor2_1 _10152_ (.A(_04393_),
    .B(net2377),
    .Y(_04444_));
 sky130_fd_sc_hs__nand2_1 _10153_ (.A(net2340),
    .B(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hs__o21ai_1 _10154_ (.A1(_04443_),
    .A2(net2339),
    .B1(_04445_),
    .Y(_04446_));
 sky130_fd_sc_hs__nand3_1 _10155_ (.A(net2328),
    .B(net2338),
    .C(_04420_),
    .Y(_04447_));
 sky130_fd_sc_hs__xnor2_1 _10156_ (.A(_04446_),
    .B(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hs__nand2_1 _10157_ (.A(_04442_),
    .B(_04448_),
    .Y(_04449_));
 sky130_fd_sc_hs__nand3_1 _10158_ (.A(net4861),
    .B(net2315),
    .C(net2327),
    .Y(_04450_));
 sky130_fd_sc_hs__nand2_2 _10159_ (.A(_04449_),
    .B(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hs__inv_1 _10160_ (.A(_04441_),
    .Y(_04452_));
 sky130_fd_sc_hs__o21ai_1 _10161_ (.A1(_04452_),
    .A2(_04437_),
    .B1(net2318),
    .Y(_04453_));
 sky130_fd_sc_hs__nand2_1 _10162_ (.A(_04453_),
    .B(net2317),
    .Y(_04454_));
 sky130_fd_sc_hs__nand2_1 _10163_ (.A(_04417_),
    .B(net2338),
    .Y(_04455_));
 sky130_fd_sc_hs__nor2_1 _10164_ (.A(net2359),
    .B(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hs__a21oi_1 _10165_ (.A1(_04456_),
    .A2(_04420_),
    .B1(net2317),
    .Y(_04457_));
 sky130_fd_sc_hs__nand2_1 _10166_ (.A(_04442_),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hs__nand2_1 _10167_ (.A(_04454_),
    .B(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hs__nor2_2 _10168_ (.A(_04451_),
    .B(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hs__nand3_2 _10169_ (.A(_04438_),
    .B(_04420_),
    .C(net2326),
    .Y(_04461_));
 sky130_fd_sc_hs__o21bai_1 _10170_ (.A1(_04452_),
    .A2(_04437_),
    .B1_N(_04420_),
    .Y(_04462_));
 sky130_fd_sc_hs__nand2_2 _10171_ (.A(_04461_),
    .B(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hs__nand2_1 _10172_ (.A(net3026),
    .B(net3024),
    .Y(_04464_));
 sky130_fd_sc_hs__xnor2_1 _10173_ (.A(net3247),
    .B(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hs__inv_1 _10174_ (.A(_04465_),
    .Y(_04466_));
 sky130_fd_sc_hs__inv_1 _10175_ (.A(net2314),
    .Y(_04467_));
 sky130_fd_sc_hs__nand3_1 _10176_ (.A(_04463_),
    .B(_04466_),
    .C(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hs__nand2_2 _10177_ (.A(_04460_),
    .B(_04468_),
    .Y(_04469_));
 sky130_fd_sc_hs__nand2_1 _10178_ (.A(_04458_),
    .B(net2316),
    .Y(_04470_));
 sky130_fd_sc_hs__nand2_1 _10179_ (.A(_04470_),
    .B(net2303),
    .Y(_04471_));
 sky130_fd_sc_hs__nand2_2 _10180_ (.A(_04469_),
    .B(_04471_),
    .Y(_04472_));
 sky130_fd_sc_hs__nand2_1 _10181_ (.A(_04472_),
    .B(_04466_),
    .Y(_04473_));
 sky130_fd_sc_hs__nand3_1 _10182_ (.A(_04469_),
    .B(_04465_),
    .C(_04471_),
    .Y(_04474_));
 sky130_fd_sc_hs__o21ai_1 _10183_ (.A1(net3158),
    .A2(net3063),
    .B1(net3024),
    .Y(_04475_));
 sky130_fd_sc_hs__xnor2_1 _10184_ (.A(net3210),
    .B(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hs__inv_1 _10185_ (.A(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hs__nand4_2 _10186_ (.A(_04473_),
    .B(_04474_),
    .C(_04477_),
    .D(net2289),
    .Y(_04478_));
 sky130_fd_sc_hs__xnor2_1 _10187_ (.A(_04420_),
    .B(net2314),
    .Y(_04479_));
 sky130_fd_sc_hs__nand2_1 _10188_ (.A(net2297),
    .B(_04479_),
    .Y(_04480_));
 sky130_fd_sc_hs__o21ai_1 _10189_ (.A1(net2314),
    .A2(net2297),
    .B1(_04480_),
    .Y(_04481_));
 sky130_fd_sc_hs__nand2_1 _10190_ (.A(net2289),
    .B(_04466_),
    .Y(_04482_));
 sky130_fd_sc_hs__xnor2_1 _10191_ (.A(_04481_),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hs__nand2_2 _10192_ (.A(_04472_),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hs__nand3_1 _10193_ (.A(_04469_),
    .B(_04471_),
    .C(_04481_),
    .Y(_04485_));
 sky130_fd_sc_hs__nand2_2 _10194_ (.A(_04484_),
    .B(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hs__nand4_1 _10195_ (.A(net2278),
    .B(net2289),
    .C(_04466_),
    .D(net2309),
    .Y(_04487_));
 sky130_fd_sc_hs__inv_1 _10196_ (.A(net2278),
    .Y(_04488_));
 sky130_fd_sc_hs__nand2_1 _10197_ (.A(net2276),
    .B(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hs__nand2_1 _10198_ (.A(_04487_),
    .B(_04489_),
    .Y(_04490_));
 sky130_fd_sc_hs__nand2_1 _10199_ (.A(_04490_),
    .B(_04472_),
    .Y(_04491_));
 sky130_fd_sc_hs__nand3_1 _10200_ (.A(_04469_),
    .B(net2278),
    .C(net2273),
    .Y(_04492_));
 sky130_fd_sc_hs__nand2_2 _10201_ (.A(_04491_),
    .B(_04492_),
    .Y(_04493_));
 sky130_fd_sc_hs__nor2_2 _10202_ (.A(_04486_),
    .B(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hs__nand2_2 _10203_ (.A(_04478_),
    .B(_04494_),
    .Y(_04495_));
 sky130_fd_sc_hs__o21ai_1 _10204_ (.A1(net2273),
    .A2(_04489_),
    .B1(net2277),
    .Y(_04496_));
 sky130_fd_sc_hs__nand2_2 _10205_ (.A(_04496_),
    .B(net2267),
    .Y(_04497_));
 sky130_fd_sc_hs__nand2_2 _10206_ (.A(_04495_),
    .B(_04497_),
    .Y(_04498_));
 sky130_fd_sc_hs__nand2_2 _10207_ (.A(_04498_),
    .B(_04477_),
    .Y(_04499_));
 sky130_fd_sc_hs__nand3_1 _10208_ (.A(_04495_),
    .B(_04476_),
    .C(_04497_),
    .Y(_04500_));
 sky130_fd_sc_hs__buf_1 place2104 (.A(_03515_),
    .X(net2104));
 sky130_fd_sc_hs__o21ai_1 _10210_ (.A1(net3120),
    .A2(net3209),
    .B1(net3024),
    .Y(_04502_));
 sky130_fd_sc_hs__xnor2_1 _10211_ (.A(net3254),
    .B(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hs__inv_1 _10212_ (.A(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hs__nand2_1 _10213_ (.A(net2254),
    .B(net2262),
    .Y(_04505_));
 sky130_fd_sc_hs__inv_1 _10214_ (.A(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hs__nand4_2 _10215_ (.A(_04499_),
    .B(_04500_),
    .C(_04504_),
    .D(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hs__nor2b_2 _10216_ (.A(_04486_),
    .B_N(_04478_),
    .Y(_04508_));
 sky130_fd_sc_hs__inv_1 _10217_ (.A(_04497_),
    .Y(_04509_));
 sky130_fd_sc_hs__nand3_1 _10218_ (.A(_04508_),
    .B(net2241),
    .C(_04509_),
    .Y(_04510_));
 sky130_fd_sc_hs__or2_1 _10219_ (.A(net2241),
    .B(_04508_),
    .X(_04511_));
 sky130_fd_sc_hs__nand2_1 _10220_ (.A(_04510_),
    .B(_04511_),
    .Y(_04512_));
 sky130_fd_sc_hs__xnor2_1 _10221_ (.A(_04465_),
    .B(net2289),
    .Y(_04513_));
 sky130_fd_sc_hs__nand2_1 _10222_ (.A(net2263),
    .B(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hs__nand3_1 _10223_ (.A(net2268),
    .B(net2289),
    .C(net2272),
    .Y(_04515_));
 sky130_fd_sc_hs__nand2_1 _10224_ (.A(_04514_),
    .B(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hs__nand3_1 _10225_ (.A(net2254),
    .B(net2262),
    .C(_04477_),
    .Y(_04517_));
 sky130_fd_sc_hs__xnor2_1 _10226_ (.A(_04516_),
    .B(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hs__nand2_1 _10227_ (.A(_04498_),
    .B(_04518_),
    .Y(_04519_));
 sky130_fd_sc_hs__nand3_1 _10228_ (.A(_04495_),
    .B(net2239),
    .C(_04497_),
    .Y(_04520_));
 sky130_fd_sc_hs__nand2_1 _10229_ (.A(_04519_),
    .B(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hs__inv_1 _10230_ (.A(net2202),
    .Y(_04522_));
 sky130_fd_sc_hs__a21o_1 _10231_ (.A1(net2203),
    .A2(_04512_),
    .B1(_04522_),
    .X(_04523_));
 sky130_fd_sc_hs__o21ai_1 _10232_ (.A1(_04509_),
    .A2(net2234),
    .B1(net2243),
    .Y(_04524_));
 sky130_fd_sc_hs__nand2_1 _10233_ (.A(_04524_),
    .B(net2242),
    .Y(_04525_));
 sky130_fd_sc_hs__nand2_1 _10234_ (.A(_04498_),
    .B(_04508_),
    .Y(_04526_));
 sky130_fd_sc_hs__and2_1 _10235_ (.A(_04525_),
    .B(_04526_),
    .X(_04527_));
 sky130_fd_sc_hs__o211ai_1 _10236_ (.A1(_04512_),
    .A2(_04527_),
    .B1(_04522_),
    .C1(_04507_),
    .Y(_04528_));
 sky130_fd_sc_hs__and2_1 _10237_ (.A(_04523_),
    .B(_04528_),
    .X(_04529_));
 sky130_fd_sc_hs__inv_2 _10238_ (.A(_04512_),
    .Y(_04530_));
 sky130_fd_sc_hs__nand2_1 _10239_ (.A(net2203),
    .B(_04522_),
    .Y(_04531_));
 sky130_fd_sc_hs__nand2_1 _10240_ (.A(_04525_),
    .B(_04526_),
    .Y(_04532_));
 sky130_fd_sc_hs__o21ai_2 _10241_ (.A1(_04530_),
    .A2(_04531_),
    .B1(net2201),
    .Y(_04533_));
 sky130_fd_sc_hs__nor2_2 _10242_ (.A(_04521_),
    .B(_04532_),
    .Y(_04534_));
 sky130_fd_sc_hs__nand2_2 _10243_ (.A(_04507_),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hs__and2_1 _10244_ (.A(_04533_),
    .B(net2193),
    .X(_04536_));
 sky130_fd_sc_hs__nand2_2 _10245_ (.A(_04535_),
    .B(_04530_),
    .Y(_04537_));
 sky130_fd_sc_hs__xnor2_1 _10246_ (.A(_04477_),
    .B(_04505_),
    .Y(_04538_));
 sky130_fd_sc_hs__nand2_1 _10247_ (.A(_04498_),
    .B(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hs__o21ai_2 _10248_ (.A1(net2240),
    .A2(net2225),
    .B1(_04539_),
    .Y(_04540_));
 sky130_fd_sc_hs__nand3_1 _10249_ (.A(net2211),
    .B(net2224),
    .C(_04504_),
    .Y(_04541_));
 sky130_fd_sc_hs__xnor2_1 _10250_ (.A(_04540_),
    .B(_04541_),
    .Y(_04542_));
 sky130_fd_sc_hs__nand2_1 _10251_ (.A(_04537_),
    .B(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hs__nand3_1 _10252_ (.A(_04535_),
    .B(_04530_),
    .C(net2200),
    .Y(_04544_));
 sky130_fd_sc_hs__nand2_1 _10253_ (.A(_04543_),
    .B(_04544_),
    .Y(_04545_));
 sky130_fd_sc_hs__inv_1 _10254_ (.A(net2161),
    .Y(_04546_));
 sky130_fd_sc_hs__nand3_1 _10255_ (.A(_04535_),
    .B(_04504_),
    .C(_04530_),
    .Y(_04547_));
 sky130_fd_sc_hs__o21ai_1 _10256_ (.A1(net2223),
    .A2(_04534_),
    .B1(_04503_),
    .Y(_04548_));
 sky130_fd_sc_hs__nand2_2 _10257_ (.A(_04547_),
    .B(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hs__nand2_1 _10258_ (.A(net3063),
    .B(net3024),
    .Y(_04550_));
 sky130_fd_sc_hs__xnor2_1 _10259_ (.A(net3202),
    .B(_04550_),
    .Y(_04551_));
 sky130_fd_sc_hs__inv_1 _10260_ (.A(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hs__nand2_1 _10261_ (.A(net2211),
    .B(net2224),
    .Y(_04553_));
 sky130_fd_sc_hs__inv_1 _10262_ (.A(_04553_),
    .Y(_04554_));
 sky130_fd_sc_hs__nand3_2 _10263_ (.A(_04554_),
    .B(_04552_),
    .C(_04549_),
    .Y(_04555_));
 sky130_fd_sc_hs__o211ai_1 _10264_ (.A1(_04529_),
    .A2(_04536_),
    .B1(_04546_),
    .C1(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hs__a21o_1 _10265_ (.A1(_04555_),
    .A2(_04536_),
    .B1(_04546_),
    .X(_04557_));
 sky130_fd_sc_hs__nand2_1 _10266_ (.A(_04556_),
    .B(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hs__nand2_1 _10267_ (.A(_04523_),
    .B(_04528_),
    .Y(_04559_));
 sky130_fd_sc_hs__nor2_2 _10268_ (.A(_04559_),
    .B(_04545_),
    .Y(_04560_));
 sky130_fd_sc_hs__nand2_2 _10269_ (.A(_04560_),
    .B(_04555_),
    .Y(_04561_));
 sky130_fd_sc_hs__nand2_2 _10270_ (.A(_04533_),
    .B(net2193),
    .Y(_04562_));
 sky130_fd_sc_hs__nand2_1 _10271_ (.A(_04561_),
    .B(_04562_),
    .Y(_04563_));
 sky130_fd_sc_hs__nand2_1 _10272_ (.A(net2185),
    .B(_04504_),
    .Y(_04564_));
 sky130_fd_sc_hs__nand3_1 _10273_ (.A(net2193),
    .B(_04503_),
    .C(net2210),
    .Y(_04565_));
 sky130_fd_sc_hs__nand2_1 _10274_ (.A(_04564_),
    .B(_04565_),
    .Y(_04566_));
 sky130_fd_sc_hs__xnor2_1 _10275_ (.A(_04504_),
    .B(_04553_),
    .Y(_04567_));
 sky130_fd_sc_hs__nand2_1 _10276_ (.A(net2185),
    .B(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hs__o21ai_1 _10277_ (.A1(_04553_),
    .A2(net2185),
    .B1(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hs__o21ai_1 _10278_ (.A1(_04551_),
    .A2(_04566_),
    .B1(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hs__nand4_1 _10279_ (.A(net2174),
    .B(net2183),
    .C(_04552_),
    .D(net2199),
    .Y(_04571_));
 sky130_fd_sc_hs__nand2_1 _10280_ (.A(_04570_),
    .B(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hs__nand2_1 _10281_ (.A(_04563_),
    .B(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hs__nand3_1 _10282_ (.A(_04561_),
    .B(_04562_),
    .C(net2158),
    .Y(_04574_));
 sky130_fd_sc_hs__nand2_2 _10283_ (.A(_04573_),
    .B(_04574_),
    .Y(_04575_));
 sky130_fd_sc_hs__nor2_4 _10284_ (.A(_04558_),
    .B(_04575_),
    .Y(_04576_));
 sky130_fd_sc_hs__nand3_1 _10285_ (.A(_04561_),
    .B(_04552_),
    .C(_04562_),
    .Y(_04577_));
 sky130_fd_sc_hs__o21ai_1 _10286_ (.A1(_04536_),
    .A2(_04560_),
    .B1(_04551_),
    .Y(_04578_));
 sky130_fd_sc_hs__nand2_2 _10287_ (.A(_04577_),
    .B(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hs__nand2_1 _10288_ (.A(net2134),
    .B(net2176),
    .Y(_04580_));
 sky130_fd_sc_hs__nand2_1 _10289_ (.A(_04576_),
    .B(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hs__nand2_1 _10290_ (.A(net3024),
    .B(net3120),
    .Y(_04582_));
 sky130_fd_sc_hs__xnor2_1 _10291_ (.A(net3201),
    .B(_04582_),
    .Y(_04583_));
 sky130_fd_sc_hs__inv_1 _10292_ (.A(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hs__nand2_1 _10293_ (.A(net2160),
    .B(_04546_),
    .Y(_04585_));
 sky130_fd_sc_hs__o21ai_1 _10294_ (.A1(_04562_),
    .A2(_04585_),
    .B1(net2184),
    .Y(_04586_));
 sky130_fd_sc_hs__and2_2 _10295_ (.A(net2152),
    .B(_04586_),
    .X(_04587_));
 sky130_fd_sc_hs__inv_1 _10296_ (.A(_04587_),
    .Y(_04588_));
 sky130_fd_sc_hs__nand3_1 _10297_ (.A(_04581_),
    .B(_04584_),
    .C(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hs__o21ai_1 _10298_ (.A1(net4901),
    .A2(_04576_),
    .B1(_04583_),
    .Y(_04590_));
 sky130_fd_sc_hs__nand2_2 _10299_ (.A(_04589_),
    .B(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hs__or2_1 _10300_ (.A(net3075),
    .B(net3112),
    .X(_04592_));
 sky130_fd_sc_hs__xnor2_1 _10301_ (.A(net3284),
    .B(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hs__inv_1 _10302_ (.A(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hs__nand3_2 _10303_ (.A(_04591_),
    .B(_04594_),
    .C(net2136),
    .Y(_04595_));
 sky130_fd_sc_hs__and2_1 _10304_ (.A(_04556_),
    .B(_04557_),
    .X(_04596_));
 sky130_fd_sc_hs__inv_1 _10305_ (.A(net2128),
    .Y(_04597_));
 sky130_fd_sc_hs__nand3_2 _10306_ (.A(_04579_),
    .B(_04584_),
    .C(net2176),
    .Y(_04598_));
 sky130_fd_sc_hs__o211ai_1 _10307_ (.A1(_04596_),
    .A2(net4900),
    .B1(_04597_),
    .C1(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hs__a21o_1 _10308_ (.A1(_04598_),
    .A2(net4900),
    .B1(_04597_),
    .X(_04600_));
 sky130_fd_sc_hs__nand2_1 _10309_ (.A(_04599_),
    .B(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hs__nand2_2 _10310_ (.A(_04598_),
    .B(_04576_),
    .Y(_04602_));
 sky130_fd_sc_hs__nand2_1 _10311_ (.A(_04602_),
    .B(_04588_),
    .Y(_04603_));
 sky130_fd_sc_hs__nand2_1 _10312_ (.A(net2144),
    .B(_04552_),
    .Y(_04604_));
 sky130_fd_sc_hs__nand2_1 _10313_ (.A(_04604_),
    .B(net2176),
    .Y(_04605_));
 sky130_fd_sc_hs__nand3_1 _10314_ (.A(net2144),
    .B(_04552_),
    .C(net2159),
    .Y(_04606_));
 sky130_fd_sc_hs__nand2_1 _10315_ (.A(_04605_),
    .B(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hs__nand2_1 _10316_ (.A(net2135),
    .B(_04584_),
    .Y(_04608_));
 sky130_fd_sc_hs__nand2_1 _10317_ (.A(_04607_),
    .B(_04608_),
    .Y(_04609_));
 sky130_fd_sc_hs__nand3_1 _10318_ (.A(net2153),
    .B(_04551_),
    .C(net2175),
    .Y(_04610_));
 sky130_fd_sc_hs__nand4_1 _10319_ (.A(_04604_),
    .B(_04610_),
    .C(_04584_),
    .D(net2159),
    .Y(_04611_));
 sky130_fd_sc_hs__nand2_1 _10320_ (.A(_04609_),
    .B(_04611_),
    .Y(_04612_));
 sky130_fd_sc_hs__nand2_1 _10321_ (.A(_04603_),
    .B(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hs__nand3_1 _10322_ (.A(_04602_),
    .B(net2126),
    .C(_04607_),
    .Y(_04614_));
 sky130_fd_sc_hs__nand2_1 _10323_ (.A(_04613_),
    .B(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hs__nor2_2 _10324_ (.A(_04601_),
    .B(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hs__nand2_2 _10325_ (.A(_04616_),
    .B(_04595_),
    .Y(_04617_));
 sky130_fd_sc_hs__nand2_1 _10326_ (.A(_04598_),
    .B(_04597_),
    .Y(_04618_));
 sky130_fd_sc_hs__o21ai_1 _10327_ (.A1(_04588_),
    .A2(_04618_),
    .B1(net2145),
    .Y(_04619_));
 sky130_fd_sc_hs__and2_2 _10328_ (.A(_04619_),
    .B(net2117),
    .X(_04620_));
 sky130_fd_sc_hs__inv_1 _10329_ (.A(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hs__nand2_2 _10330_ (.A(_04617_),
    .B(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hs__nand2_2 _10331_ (.A(_04622_),
    .B(_04594_),
    .Y(_04623_));
 sky130_fd_sc_hs__nand3_1 _10332_ (.A(_04617_),
    .B(_04593_),
    .C(_04621_),
    .Y(_04624_));
 sky130_fd_sc_hs__or2_1 _10333_ (.A(net3163),
    .B(net3075),
    .X(_04625_));
 sky130_fd_sc_hs__xnor2_1 _10334_ (.A(net3250),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hs__inv_1 _10335_ (.A(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hs__nand4_1 _10336_ (.A(_04623_),
    .B(_04624_),
    .C(_04627_),
    .D(net2099),
    .Y(_04628_));
 sky130_fd_sc_hs__and2_1 _10337_ (.A(_04599_),
    .B(_04600_),
    .X(_04629_));
 sky130_fd_sc_hs__inv_1 _10338_ (.A(_04615_),
    .Y(_04630_));
 sky130_fd_sc_hs__o211ai_1 _10339_ (.A1(_04629_),
    .A2(_04620_),
    .B1(_04630_),
    .C1(_04595_),
    .Y(_04631_));
 sky130_fd_sc_hs__a21o_1 _10340_ (.A1(_04595_),
    .A2(_04620_),
    .B1(_04630_),
    .X(_04632_));
 sky130_fd_sc_hs__nand2_1 _10341_ (.A(_04631_),
    .B(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hs__xnor2_1 _10342_ (.A(_04583_),
    .B(net2136),
    .Y(_04634_));
 sky130_fd_sc_hs__nand2_1 _10343_ (.A(net2109),
    .B(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hs__nand3_1 _10344_ (.A(net2118),
    .B(net2136),
    .C(net2127),
    .Y(_04636_));
 sky130_fd_sc_hs__nand2_1 _10345_ (.A(_04635_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hs__nand2_1 _10346_ (.A(net2098),
    .B(_04594_),
    .Y(_04638_));
 sky130_fd_sc_hs__xnor2_1 _10347_ (.A(_04637_),
    .B(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hs__nand2_1 _10348_ (.A(_04622_),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hs__nand3_1 _10349_ (.A(_04617_),
    .B(net2089),
    .C(_04621_),
    .Y(_04641_));
 sky130_fd_sc_hs__nand2_1 _10350_ (.A(_04640_),
    .B(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hs__nor2_1 _10351_ (.A(_04633_),
    .B(_04642_),
    .Y(_04643_));
 sky130_fd_sc_hs__nand2_2 _10352_ (.A(_04628_),
    .B(_04643_),
    .Y(_04644_));
 sky130_fd_sc_hs__nand2_1 _10353_ (.A(net2079),
    .B(net2110),
    .Y(_04645_));
 sky130_fd_sc_hs__nand2_4 _10354_ (.A(_04645_),
    .B(net2080),
    .Y(_04646_));
 sky130_fd_sc_hs__nand2_2 _10355_ (.A(_04644_),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hs__nand3_1 _10356_ (.A(_04623_),
    .B(_04624_),
    .C(net2099),
    .Y(_04648_));
 sky130_fd_sc_hs__nor2_1 _10357_ (.A(_04626_),
    .B(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hs__nor2_1 _10358_ (.A(net2054),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hs__nand2_1 _10359_ (.A(_04647_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hs__inv_1 _10360_ (.A(net2071),
    .Y(_04652_));
 sky130_fd_sc_hs__nand2_1 _10361_ (.A(_04651_),
    .B(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hs__inv_1 _10362_ (.A(net2063),
    .Y(_04654_));
 sky130_fd_sc_hs__nand3_1 _10363_ (.A(net2044),
    .B(net2071),
    .C(_04654_),
    .Y(_04655_));
 sky130_fd_sc_hs__nand2_1 _10364_ (.A(_04653_),
    .B(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hs__o21ai_1 _10365_ (.A1(_04646_),
    .A2(_04649_),
    .B1(net2054),
    .Y(_04657_));
 sky130_fd_sc_hs__nand2_1 _10366_ (.A(_04651_),
    .B(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hs__inv_1 _10367_ (.A(net2099),
    .Y(_04659_));
 sky130_fd_sc_hs__nand2_1 _10368_ (.A(_04623_),
    .B(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hs__nand3_1 _10369_ (.A(_04622_),
    .B(_04594_),
    .C(net2099),
    .Y(_04661_));
 sky130_fd_sc_hs__and2_1 _10370_ (.A(_04660_),
    .B(_04661_),
    .X(_04662_));
 sky130_fd_sc_hs__and2_2 _10371_ (.A(_04623_),
    .B(_04624_),
    .X(_04663_));
 sky130_fd_sc_hs__nand2_1 _10372_ (.A(_04663_),
    .B(_04627_),
    .Y(_04664_));
 sky130_fd_sc_hs__nand2_1 _10373_ (.A(_04662_),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hs__nand2_1 _10374_ (.A(_04623_),
    .B(_04624_),
    .Y(_04666_));
 sky130_fd_sc_hs__nor2_1 _10375_ (.A(_04626_),
    .B(_04666_),
    .Y(_04667_));
 sky130_fd_sc_hs__nand2_1 _10376_ (.A(_04660_),
    .B(_04661_),
    .Y(_04668_));
 sky130_fd_sc_hs__nand2_1 _10377_ (.A(_04667_),
    .B(_04668_),
    .Y(_04669_));
 sky130_fd_sc_hs__nand2_1 _10378_ (.A(_04665_),
    .B(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hs__nand2_1 _10379_ (.A(_04647_),
    .B(_04670_),
    .Y(_04671_));
 sky130_fd_sc_hs__nand3_1 _10380_ (.A(_04644_),
    .B(_04662_),
    .C(_04646_),
    .Y(_04672_));
 sky130_fd_sc_hs__nand2_2 _10381_ (.A(_04671_),
    .B(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hs__nor2_2 _10382_ (.A(_04658_),
    .B(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hs__nand2_1 _10383_ (.A(_04647_),
    .B(_04627_),
    .Y(_04675_));
 sky130_fd_sc_hs__nand3_1 _10384_ (.A(_04644_),
    .B(_04626_),
    .C(_04646_),
    .Y(_04676_));
 sky130_fd_sc_hs__nand2_1 _10385_ (.A(net3024),
    .B(net3156),
    .Y(_04677_));
 sky130_fd_sc_hs__xnor2_1 _10386_ (.A(net3285),
    .B(_04677_),
    .Y(_04678_));
 sky130_fd_sc_hs__nand4_2 _10387_ (.A(_04675_),
    .B(_04676_),
    .C(_04678_),
    .D(net2053),
    .Y(_04679_));
 sky130_fd_sc_hs__o211ai_1 _10388_ (.A1(net2003),
    .A2(net2002),
    .B1(net2008),
    .C1(net2007),
    .Y(_04680_));
 sky130_fd_sc_hs__o21ai_1 _10389_ (.A1(net2003),
    .A2(net2002),
    .B1(net2007),
    .Y(_04681_));
 sky130_fd_sc_hs__inv_1 _10390_ (.A(_04673_),
    .Y(_04682_));
 sky130_fd_sc_hs__nand2_1 _10391_ (.A(_04681_),
    .B(net2001),
    .Y(_04683_));
 sky130_fd_sc_hs__nand2_1 _10392_ (.A(_04680_),
    .B(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hs__inv_1 _10393_ (.A(_04656_),
    .Y(_04685_));
 sky130_fd_sc_hs__nand2_1 _10394_ (.A(_04679_),
    .B(_04682_),
    .Y(_04686_));
 sky130_fd_sc_hs__o21ai_1 _10395_ (.A1(_04685_),
    .A2(_04686_),
    .B1(net2009),
    .Y(_04687_));
 sky130_fd_sc_hs__nand2_2 _10396_ (.A(_04679_),
    .B(_04674_),
    .Y(_04688_));
 sky130_fd_sc_hs__and2_2 _10397_ (.A(_04687_),
    .B(net1994),
    .X(_04689_));
 sky130_fd_sc_hs__nand2_2 _10398_ (.A(_04688_),
    .B(_04685_),
    .Y(_04690_));
 sky130_fd_sc_hs__a21oi_1 _10399_ (.A1(net2045),
    .A2(net2064),
    .B1(net2050),
    .Y(_04691_));
 sky130_fd_sc_hs__a21oi_1 _10400_ (.A1(net2035),
    .A2(_04627_),
    .B1(net2053),
    .Y(_04692_));
 sky130_fd_sc_hs__nor2_1 _10401_ (.A(_04691_),
    .B(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hs__and2_2 _10402_ (.A(net2021),
    .B(net2034),
    .X(_04694_));
 sky130_fd_sc_hs__nand2_1 _10403_ (.A(_04694_),
    .B(_04678_),
    .Y(_04695_));
 sky130_fd_sc_hs__nand2_1 _10404_ (.A(_04693_),
    .B(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hs__nand4_1 _10405_ (.A(net2021),
    .B(net2034),
    .C(_04678_),
    .D(net2052),
    .Y(_04697_));
 sky130_fd_sc_hs__nand2_1 _10406_ (.A(_04696_),
    .B(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hs__nand2_1 _10407_ (.A(_04690_),
    .B(_04698_),
    .Y(_04699_));
 sky130_fd_sc_hs__nand3_1 _10408_ (.A(net1995),
    .B(net1998),
    .C(_04693_),
    .Y(_04700_));
 sky130_fd_sc_hs__and2_2 _10409_ (.A(_04699_),
    .B(_04700_),
    .X(_04701_));
 sky130_fd_sc_hs__nand2_1 _10410_ (.A(_04690_),
    .B(_04678_),
    .Y(_04702_));
 sky130_fd_sc_hs__inv_1 _10411_ (.A(_04678_),
    .Y(_04703_));
 sky130_fd_sc_hs__nand3_1 _10412_ (.A(net1996),
    .B(_04703_),
    .C(net1998),
    .Y(_04704_));
 sky130_fd_sc_hs__nor2_1 _10413_ (.A(net3252),
    .B(net3075),
    .Y(_04705_));
 sky130_fd_sc_hs__xnor2_1 _10414_ (.A(net3325),
    .B(_04705_),
    .Y(_04706_));
 sky130_fd_sc_hs__nand4_1 _10415_ (.A(_04702_),
    .B(_04704_),
    .C(_04706_),
    .D(net2006),
    .Y(_04707_));
 sky130_fd_sc_hs__o211ai_1 _10416_ (.A1(net1978),
    .A2(_04689_),
    .B1(net1966),
    .C1(net1965),
    .Y(_04708_));
 sky130_fd_sc_hs__a21o_1 _10417_ (.A1(_04707_),
    .A2(_04689_),
    .B1(net1966),
    .X(_04709_));
 sky130_fd_sc_hs__nand2_1 _10418_ (.A(_04708_),
    .B(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hs__nand2_1 _10419_ (.A(_04699_),
    .B(_04700_),
    .Y(_04711_));
 sky130_fd_sc_hs__nand4_1 _10420_ (.A(_04694_),
    .B(net2008),
    .C(_04678_),
    .D(net2053),
    .Y(_04712_));
 sky130_fd_sc_hs__nand2_1 _10421_ (.A(_04712_),
    .B(_04686_),
    .Y(_04713_));
 sky130_fd_sc_hs__nand2_1 _10422_ (.A(_04713_),
    .B(_04690_),
    .Y(_04714_));
 sky130_fd_sc_hs__nand3_1 _10423_ (.A(_04688_),
    .B(_04685_),
    .C(net2008),
    .Y(_04715_));
 sky130_fd_sc_hs__nand2_1 _10424_ (.A(_04714_),
    .B(_04715_),
    .Y(_04716_));
 sky130_fd_sc_hs__nor2_2 _10425_ (.A(_04711_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hs__nand2_2 _10426_ (.A(_04707_),
    .B(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hs__inv_1 _10427_ (.A(_04689_),
    .Y(_04719_));
 sky130_fd_sc_hs__nand2_2 _10428_ (.A(_04718_),
    .B(_04719_),
    .Y(_04720_));
 sky130_fd_sc_hs__inv_1 _10429_ (.A(_04706_),
    .Y(_04721_));
 sky130_fd_sc_hs__nand2_1 _10430_ (.A(_04702_),
    .B(net1985),
    .Y(_04722_));
 sky130_fd_sc_hs__nor2_1 _10431_ (.A(_04721_),
    .B(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hs__xnor2_1 _10432_ (.A(_04703_),
    .B(net2006),
    .Y(_04724_));
 sky130_fd_sc_hs__nand2_1 _10433_ (.A(net1986),
    .B(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hs__nand3_1 _10434_ (.A(net1997),
    .B(net1998),
    .C(net2006),
    .Y(_04726_));
 sky130_fd_sc_hs__nand2_1 _10435_ (.A(_04725_),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hs__inv_1 _10436_ (.A(_04727_),
    .Y(_04728_));
 sky130_fd_sc_hs__nand2_1 _10437_ (.A(_04723_),
    .B(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hs__o21ai_1 _10438_ (.A1(_04721_),
    .A2(_04722_),
    .B1(_04727_),
    .Y(_04730_));
 sky130_fd_sc_hs__nand2_1 _10439_ (.A(_04729_),
    .B(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hs__nand2_1 _10440_ (.A(_04720_),
    .B(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hs__nand3_1 _10441_ (.A(_04718_),
    .B(_04719_),
    .C(_04727_),
    .Y(_04733_));
 sky130_fd_sc_hs__nand2_2 _10442_ (.A(_04732_),
    .B(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hs__nor2_2 _10443_ (.A(_04710_),
    .B(_04734_),
    .Y(_04735_));
 sky130_fd_sc_hs__nand3_1 _10444_ (.A(_04702_),
    .B(_04704_),
    .C(net2006),
    .Y(_04736_));
 sky130_fd_sc_hs__nand3_1 _10445_ (.A(_04736_),
    .B(_04701_),
    .C(_04684_),
    .Y(_04737_));
 sky130_fd_sc_hs__nand3_1 _10446_ (.A(_04737_),
    .B(_04706_),
    .C(_04719_),
    .Y(_04738_));
 sky130_fd_sc_hs__o21ai_2 _10447_ (.A1(_04689_),
    .A2(_04717_),
    .B1(_04721_),
    .Y(_04739_));
 sky130_fd_sc_hs__nand2_1 _10448_ (.A(_04738_),
    .B(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hs__nor2_1 _10449_ (.A(net3283),
    .B(net3075),
    .Y(_04741_));
 sky130_fd_sc_hs__xnor2_1 _10450_ (.A(net3286),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hs__inv_1 _10451_ (.A(net1963),
    .Y(_04743_));
 sky130_fd_sc_hs__nand3_1 _10452_ (.A(_04740_),
    .B(_04742_),
    .C(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hs__nand2_2 _10453_ (.A(_04735_),
    .B(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hs__nand2_1 _10454_ (.A(_04708_),
    .B(net1964),
    .Y(_04746_));
 sky130_fd_sc_hs__nand2_1 _10455_ (.A(_04746_),
    .B(net1955),
    .Y(_04747_));
 sky130_fd_sc_hs__nand2_2 _10456_ (.A(_04745_),
    .B(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hs__nand2_2 _10457_ (.A(_04748_),
    .B(_04742_),
    .Y(_04749_));
 sky130_fd_sc_hs__nand3b_1 _10458_ (.A_N(_04742_),
    .B(_04745_),
    .C(_04747_),
    .Y(_04750_));
 sky130_fd_sc_hs__nand3_1 _10459_ (.A(_04749_),
    .B(_04750_),
    .C(net1947),
    .Y(_04751_));
 sky130_fd_sc_hs__a21boi_1 _10460_ (.A1(net1954),
    .A2(net1953),
    .B1_N(_04743_),
    .Y(_04752_));
 sky130_fd_sc_hs__nand3_1 _10461_ (.A(_04752_),
    .B(_04742_),
    .C(net1923),
    .Y(_04753_));
 sky130_fd_sc_hs__inv_2 _10462_ (.A(_04734_),
    .Y(_04754_));
 sky130_fd_sc_hs__nand2_1 _10463_ (.A(_04754_),
    .B(net1936),
    .Y(_04755_));
 sky130_fd_sc_hs__nand2_1 _10464_ (.A(_04753_),
    .B(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hs__nand2_1 _10465_ (.A(_04756_),
    .B(_04748_),
    .Y(_04757_));
 sky130_fd_sc_hs__nand3_1 _10466_ (.A(_04745_),
    .B(_04747_),
    .C(net1923),
    .Y(_04758_));
 sky130_fd_sc_hs__nand2_2 _10467_ (.A(_04757_),
    .B(_04758_),
    .Y(_04759_));
 sky130_fd_sc_hs__nand2_1 _10468_ (.A(_04740_),
    .B(_04742_),
    .Y(_04760_));
 sky130_fd_sc_hs__xnor2_1 _10469_ (.A(_04706_),
    .B(_04722_),
    .Y(_04761_));
 sky130_fd_sc_hs__nand2_1 _10470_ (.A(_04720_),
    .B(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hs__o21ai_1 _10471_ (.A1(net1963),
    .A2(_04720_),
    .B1(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hs__or2_1 _10472_ (.A(_04760_),
    .B(_04763_),
    .X(_04764_));
 sky130_fd_sc_hs__nand2_1 _10473_ (.A(_04763_),
    .B(net1935),
    .Y(_04765_));
 sky130_fd_sc_hs__nand2_1 _10474_ (.A(_04764_),
    .B(_04765_),
    .Y(_04766_));
 sky130_fd_sc_hs__nand2_1 _10475_ (.A(_04748_),
    .B(_04766_),
    .Y(_04767_));
 sky130_fd_sc_hs__nand3_1 _10476_ (.A(_04745_),
    .B(_04763_),
    .C(_04747_),
    .Y(_04768_));
 sky130_fd_sc_hs__nand2_1 _10477_ (.A(_04767_),
    .B(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hs__nand2_1 _10478_ (.A(_04759_),
    .B(_04769_),
    .Y(_04770_));
 sky130_fd_sc_hs__nor3_2 _10479_ (.A(_03928_),
    .B(_04751_),
    .C(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hs__a21oi_1 _10480_ (.A1(_04747_),
    .A2(net1956),
    .B1(net1917),
    .Y(_04772_));
 sky130_fd_sc_hs__xor2_2 _10481_ (.A(net1956),
    .B(_04772_),
    .X(_04773_));
 sky130_fd_sc_hs__a21oi_2 _10482_ (.A1(net1871),
    .A2(net1896),
    .B1(net3075),
    .Y(_04774_));
 sky130_fd_sc_hs__nor2_8 _10483_ (.A(net1845),
    .B(_04774_),
    .Y(_04775_));
 sky130_fd_sc_hs__buf_1 place2103 (.A(_03521_),
    .X(net2103));
 sky130_fd_sc_hs__a211oi_2 _10485_ (.A1(net4962),
    .A2(net3605),
    .B1(net3782),
    .C1(net4972),
    .Y(_00492_));
 sky130_fd_sc_hs__nand2_1 _10486_ (.A(net1896),
    .B(net1887),
    .Y(_04777_));
 sky130_fd_sc_hs__inv_1 _10487_ (.A(net3329),
    .Y(_04778_));
 sky130_fd_sc_hs__nand2_1 _10488_ (.A(net3024),
    .B(net3603),
    .Y(_04779_));
 sky130_fd_sc_hs__o2111ai_1 _10489_ (.A1(net3024),
    .A2(_04778_),
    .B1(net3442),
    .C1(_04779_),
    .D1(_03927_),
    .Y(_04780_));
 sky130_fd_sc_hs__nand2_1 _10490_ (.A(net1898),
    .B(net1908),
    .Y(_04781_));
 sky130_fd_sc_hs__nor2_2 _10491_ (.A(_04780_),
    .B(_04781_),
    .Y(_04782_));
 sky130_fd_sc_hs__nand3_2 _10492_ (.A(_04782_),
    .B(net1947),
    .C(net1886),
    .Y(_04783_));
 sky130_fd_sc_hs__o21a_4 _10493_ (.A1(_04777_),
    .A2(_04783_),
    .B1(net3024),
    .X(_04784_));
 sky130_fd_sc_hs__o21ai_1 _10494_ (.A1(net1845),
    .A2(_04784_),
    .B1(net3784),
    .Y(_04785_));
 sky130_fd_sc_hs__a21oi_1 _10495_ (.A1(net3577),
    .A2(net4973),
    .B1(_04785_),
    .Y(_00493_));
 sky130_fd_sc_hs__a211oi_4 _10496_ (.A1(net4962),
    .A2(net3581),
    .B1(net3782),
    .C1(net4972),
    .Y(_00494_));
 sky130_fd_sc_hs__buf_1 place2105 (.A(net3797),
    .X(net2105));
 sky130_fd_sc_hs__nor2_8 _10498_ (.A(net1845),
    .B(_04784_),
    .Y(_04787_));
 sky130_fd_sc_hs__a211oi_4 _10499_ (.A1(net4973),
    .A2(net3582),
    .B1(net3782),
    .C1(net4961),
    .Y(_00495_));
 sky130_fd_sc_hs__a211oi_4 _10500_ (.A1(net4962),
    .A2(net3576),
    .B1(net3782),
    .C1(net4972),
    .Y(_00496_));
 sky130_fd_sc_hs__a211oi_2 _10501_ (.A1(net4973),
    .A2(net3575),
    .B1(net3782),
    .C1(net4961),
    .Y(_00497_));
 sky130_fd_sc_hs__a211oi_2 _10502_ (.A1(net4962),
    .A2(net3574),
    .B1(net3782),
    .C1(net4972),
    .Y(_00498_));
 sky130_fd_sc_hs__a211oi_2 _10503_ (.A1(net1847),
    .A2(net3591),
    .B1(net3782),
    .C1(net4961),
    .Y(_00499_));
 sky130_fd_sc_hs__a211oi_4 _10504_ (.A1(net3592),
    .A2(net1847),
    .B1(net3782),
    .C1(net3788),
    .Y(_00500_));
 sky130_fd_sc_hs__a211oi_4 _10505_ (.A1(net4962),
    .A2(net3586),
    .B1(net3782),
    .C1(net4958),
    .Y(_00501_));
 sky130_fd_sc_hs__o21ai_4 _10506_ (.A1(net3499),
    .A2(net1846),
    .B1(net3784),
    .Y(_04788_));
 sky130_fd_sc_hs__a21oi_2 _10507_ (.A1(net3602),
    .A2(net1846),
    .B1(_04788_),
    .Y(_00502_));
 sky130_fd_sc_hs__a211oi_4 _10508_ (.A1(net4962),
    .A2(net3587),
    .B1(net3782),
    .C1(net4972),
    .Y(_00503_));
 sky130_fd_sc_hs__a211oi_4 _10509_ (.A1(net4973),
    .A2(net3583),
    .B1(net3782),
    .C1(net4961),
    .Y(_00504_));
 sky130_fd_sc_hs__a211oi_4 _10510_ (.A1(net3584),
    .A2(net1847),
    .B1(net3782),
    .C1(net3788),
    .Y(_00505_));
 sky130_fd_sc_hs__bufbuf_8 place2102 (.A(_03523_),
    .X(net2102));
 sky130_fd_sc_hs__a211oi_4 _10512_ (.A1(net1847),
    .A2(net3593),
    .B1(net3783),
    .C1(net4958),
    .Y(_00506_));
 sky130_fd_sc_hs__a211oi_2 _10513_ (.A1(net3594),
    .A2(net1847),
    .B1(net3783),
    .C1(net3788),
    .Y(_00507_));
 sky130_fd_sc_hs__a211oi_2 _10514_ (.A1(net1847),
    .A2(net3595),
    .B1(net3783),
    .C1(net4958),
    .Y(_00508_));
 sky130_fd_sc_hs__a211oi_4 _10515_ (.A1(net3596),
    .A2(net1847),
    .B1(net3783),
    .C1(net3788),
    .Y(_00509_));
 sky130_fd_sc_hs__a211oi_2 _10516_ (.A1(net1847),
    .A2(net3597),
    .B1(net3783),
    .C1(net4958),
    .Y(_00510_));
 sky130_fd_sc_hs__a211oi_2 _10517_ (.A1(_03888_),
    .A2(net1847),
    .B1(net3783),
    .C1(net3788),
    .Y(_00511_));
 sky130_fd_sc_hs__a211oi_4 _10518_ (.A1(net1847),
    .A2(net3599),
    .B1(net3783),
    .C1(net4958),
    .Y(_00512_));
 sky130_fd_sc_hs__clkinv_1 _10519_ (.A(\u_hamming_window.rd_en_o ),
    .Y(_04790_));
 sky130_fd_sc_hs__nand2_2 _10520_ (.A(net4903),
    .B(\u_window_buffer.next_state_is_valid_to_read ),
    .Y(_04791_));
 sky130_fd_sc_hs__nor2_4 _10521_ (.A(_04791_),
    .B(_04790_),
    .Y(_04792_));
 sky130_fd_sc_hs__buf_1 place2100 (.A(_03542_),
    .X(net2100));
 sky130_fd_sc_hs__o21ai_4 _10523_ (.A1(net3723),
    .A2(net1842),
    .B1(net3784),
    .Y(_04794_));
 sky130_fd_sc_hs__a21oi_4 _10524_ (.A1(net4974),
    .A2(_04778_),
    .B1(_04794_),
    .Y(_00513_));
 sky130_fd_sc_hs__a211oi_4 _10525_ (.A1(net3601),
    .A2(net1847),
    .B1(net3783),
    .C1(net3788),
    .Y(_00514_));
 sky130_fd_sc_hs__nor2_2 _10526_ (.A(net3721),
    .B(net1842),
    .Y(_04795_));
 sky130_fd_sc_hs__nor3_2 _10527_ (.A(net3782),
    .B(_04795_),
    .C(net4961),
    .Y(_00515_));
 sky130_fd_sc_hs__o21ai_1 _10528_ (.A1(net3603),
    .A2(net3378),
    .B1(net3024),
    .Y(_04796_));
 sky130_fd_sc_hs__xnor2_1 _10529_ (.A(_04796_),
    .B(_03927_),
    .Y(_04797_));
 sky130_fd_sc_hs__o21ai_4 _10530_ (.A1(net3720),
    .A2(net1842),
    .B1(net3784),
    .Y(_04798_));
 sky130_fd_sc_hs__a21oi_2 _10531_ (.A1(net4974),
    .A2(_04797_),
    .B1(_04798_),
    .Y(_00516_));
 sky130_fd_sc_hs__a21oi_1 _10532_ (.A1(_03927_),
    .A2(net3377),
    .B1(net3075),
    .Y(_04799_));
 sky130_fd_sc_hs__xnor2_1 _10533_ (.A(_04799_),
    .B(net1885),
    .Y(_04800_));
 sky130_fd_sc_hs__nor2_4 _10534_ (.A(net3719),
    .B(net1842),
    .Y(_04801_));
 sky130_fd_sc_hs__a211oi_4 _10535_ (.A1(net4974),
    .A2(_04800_),
    .B1(net3782),
    .C1(_04801_),
    .Y(_00517_));
 sky130_fd_sc_hs__inv_1 _10536_ (.A(net1947),
    .Y(_04802_));
 sky130_fd_sc_hs__xnor2_1 _10537_ (.A(_04802_),
    .B(net1898),
    .Y(_04803_));
 sky130_fd_sc_hs__nor2_1 _10538_ (.A(net3075),
    .B(net1879),
    .Y(_04804_));
 sky130_fd_sc_hs__xnor2_1 _10539_ (.A(_04803_),
    .B(_04804_),
    .Y(_04805_));
 sky130_fd_sc_hs__o21ai_4 _10540_ (.A1(net3718),
    .A2(net1842),
    .B1(net3784),
    .Y(_04806_));
 sky130_fd_sc_hs__a21oi_2 _10541_ (.A1(net4974),
    .A2(_04805_),
    .B1(_04806_),
    .Y(_00518_));
 sky130_fd_sc_hs__o21ai_1 _10542_ (.A1(_03928_),
    .A2(net1888),
    .B1(net3024),
    .Y(_04807_));
 sky130_fd_sc_hs__xnor2_1 _10543_ (.A(net1886),
    .B(_04807_),
    .Y(_04808_));
 sky130_fd_sc_hs__o21ai_4 _10544_ (.A1(net3717),
    .A2(net1842),
    .B1(net3784),
    .Y(_04809_));
 sky130_fd_sc_hs__a21oi_1 _10545_ (.A1(net4974),
    .A2(_04808_),
    .B1(_04809_),
    .Y(_00519_));
 sky130_fd_sc_hs__nand2_1 _10546_ (.A(_04783_),
    .B(net3024),
    .Y(_04810_));
 sky130_fd_sc_hs__xnor2_1 _10547_ (.A(net1887),
    .B(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hs__o21ai_4 _10548_ (.A1(net3716),
    .A2(net1842),
    .B1(net3784),
    .Y(_04812_));
 sky130_fd_sc_hs__a21oi_1 _10549_ (.A1(net4974),
    .A2(_04811_),
    .B1(_04812_),
    .Y(_00520_));
 sky130_fd_sc_hs__nor2_1 _10550_ (.A(net3075),
    .B(net1871),
    .Y(_04813_));
 sky130_fd_sc_hs__xor2_1 _10551_ (.A(net1897),
    .B(_04813_),
    .X(_04814_));
 sky130_fd_sc_hs__o21ai_4 _10552_ (.A1(net3715),
    .A2(net1842),
    .B1(net3784),
    .Y(_04815_));
 sky130_fd_sc_hs__a21oi_2 _10553_ (.A1(net4974),
    .A2(_04814_),
    .B1(_04815_),
    .Y(_00521_));
 sky130_fd_sc_hs__a21oi_2 _10554_ (.A1(net3589),
    .A2(net4973),
    .B1(_04785_),
    .Y(_00522_));
 sky130_fd_sc_hs__nor2_1 _10555_ (.A(net3782),
    .B(_00658_),
    .Y(_00523_));
 sky130_fd_sc_hs__buf_1 place2101 (.A(_03536_),
    .X(net2101));
 sky130_fd_sc_hs__inv_2 _10557_ (.A(\u_window_buffer.write_ptr[0] ),
    .Y(_04817_));
 sky130_fd_sc_hs__o21ai_1 _10558_ (.A1(net3674),
    .A2(net3571),
    .B1(net3785),
    .Y(_04818_));
 sky130_fd_sc_hs__a21oi_1 _10559_ (.A1(net3674),
    .A2(net3571),
    .B1(_04818_),
    .Y(_00524_));
 sky130_fd_sc_hs__nor2_1 _10560_ (.A(net3652),
    .B(net3653),
    .Y(_04819_));
 sky130_fd_sc_hs__nor2_1 _10561_ (.A(net3661),
    .B(_02019_),
    .Y(_04820_));
 sky130_fd_sc_hs__nand2_1 _10562_ (.A(net3430),
    .B(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hs__nor2_1 _10563_ (.A(_02087_),
    .B(_02084_),
    .Y(_04822_));
 sky130_fd_sc_hs__nand3_1 _10564_ (.A(_04822_),
    .B(net3712),
    .C(net3711),
    .Y(_04823_));
 sky130_fd_sc_hs__inv_2 _10565_ (.A(\u_window_buffer.write_ptr[5] ),
    .Y(_04824_));
 sky130_fd_sc_hs__inv_2 _10566_ (.A(\u_window_buffer.write_ptr[2] ),
    .Y(_04825_));
 sky130_fd_sc_hs__inv_2 _10567_ (.A(_00228_),
    .Y(_04826_));
 sky130_fd_sc_hs__nor2_4 _10568_ (.A(_04825_),
    .B(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hs__nand2_2 _10569_ (.A(_04827_),
    .B(\u_window_buffer.write_ptr[3] ),
    .Y(_04828_));
 sky130_fd_sc_hs__nor3_4 _10570_ (.A(_02067_),
    .B(_04828_),
    .C(net3569),
    .Y(_04829_));
 sky130_fd_sc_hs__inv_1 _10571_ (.A(\u_window_buffer.write_ptr[6] ),
    .Y(_04830_));
 sky130_fd_sc_hs__nand2_1 _10572_ (.A(\u_window_buffer.write_ptr[8] ),
    .B(\u_window_buffer.write_ptr[9] ),
    .Y(_04831_));
 sky130_fd_sc_hs__nor3_1 _10573_ (.A(net3567),
    .B(_02048_),
    .C(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hs__nand2_2 _10574_ (.A(_04832_),
    .B(_04829_),
    .Y(_04833_));
 sky130_fd_sc_hs__nor2_4 _10575_ (.A(net3246),
    .B(_04823_),
    .Y(_04834_));
 sky130_fd_sc_hs__nor2_1 _10576_ (.A(_02077_),
    .B(_02073_),
    .Y(_04835_));
 sky130_fd_sc_hs__nor2_1 _10577_ (.A(_02028_),
    .B(net3657),
    .Y(_04836_));
 sky130_fd_sc_hs__nand3_2 _10578_ (.A(net3427),
    .B(_04834_),
    .C(_04836_),
    .Y(_04837_));
 sky130_fd_sc_hs__nor2_4 _10579_ (.A(_04837_),
    .B(_04821_),
    .Y(_04838_));
 sky130_fd_sc_hs__nand2_1 _10580_ (.A(\u_window_buffer.write_ptr[22] ),
    .B(\u_window_buffer.write_ptr[23] ),
    .Y(_04839_));
 sky130_fd_sc_hs__nor3_1 _10581_ (.A(_01980_),
    .B(_01976_),
    .C(_04839_),
    .Y(_04840_));
 sky130_fd_sc_hs__nand2_2 _10582_ (.A(_04838_),
    .B(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hs__xnor2_2 _10583_ (.A(_04841_),
    .B(net3667),
    .Y(_04842_));
 sky130_fd_sc_hs__nand2_1 _10584_ (.A(\u_window_buffer.write_ptr[28] ),
    .B(\u_window_buffer.write_ptr[29] ),
    .Y(_04843_));
 sky130_fd_sc_hs__nor3_1 _10585_ (.A(_01950_),
    .B(_01989_),
    .C(_04843_),
    .Y(_04844_));
 sky130_fd_sc_hs__nand2_1 _10586_ (.A(\u_window_buffer.write_ptr[23] ),
    .B(\u_window_buffer.write_ptr[24] ),
    .Y(_04845_));
 sky130_fd_sc_hs__nor3_1 _10587_ (.A(_01976_),
    .B(_01965_),
    .C(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hs__nand2_1 _10588_ (.A(_04844_),
    .B(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hs__nor2_1 _10589_ (.A(_02034_),
    .B(_02015_),
    .Y(_04848_));
 sky130_fd_sc_hs__nand3_1 _10590_ (.A(net3426),
    .B(net3699),
    .C(\u_window_buffer.write_ptr[22] ),
    .Y(_04849_));
 sky130_fd_sc_hs__nor2_1 _10591_ (.A(_02104_),
    .B(_02111_),
    .Y(_04850_));
 sky130_fd_sc_hs__inv_1 _10592_ (.A(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hs__nor2_1 _10593_ (.A(_02048_),
    .B(_02095_),
    .Y(_04852_));
 sky130_fd_sc_hs__inv_2 _10594_ (.A(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hs__nor2_1 _10595_ (.A(_04824_),
    .B(_04830_),
    .Y(_04854_));
 sky130_fd_sc_hs__inv_1 _10596_ (.A(_04854_),
    .Y(_04855_));
 sky130_fd_sc_hs__nand2_1 _10597_ (.A(\u_window_buffer.write_ptr[1] ),
    .B(\u_window_buffer.write_ptr[2] ),
    .Y(_04856_));
 sky130_fd_sc_hs__nor2_2 _10598_ (.A(_04817_),
    .B(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hs__nand3_2 _10599_ (.A(_04857_),
    .B(\u_window_buffer.write_ptr[3] ),
    .C(\u_window_buffer.write_ptr[4] ),
    .Y(_04858_));
 sky130_fd_sc_hs__or2_2 _10600_ (.A(_04855_),
    .B(_04858_),
    .X(_04859_));
 sky130_fd_sc_hs__nor3_2 _10601_ (.A(_04851_),
    .B(_04853_),
    .C(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hs__nor2_1 _10602_ (.A(_02025_),
    .B(_02038_),
    .Y(_04861_));
 sky130_fd_sc_hs__nor2_1 _10603_ (.A(net3635),
    .B(_02087_),
    .Y(_04862_));
 sky130_fd_sc_hs__inv_1 _10604_ (.A(_04862_),
    .Y(_04863_));
 sky130_fd_sc_hs__nor2_1 _10605_ (.A(_02084_),
    .B(_02077_),
    .Y(_04864_));
 sky130_fd_sc_hs__nand3_1 _10606_ (.A(_04864_),
    .B(\u_window_buffer.write_ptr[15] ),
    .C(\u_window_buffer.write_ptr[16] ),
    .Y(_04865_));
 sky130_fd_sc_hs__nor2_1 _10607_ (.A(net3369),
    .B(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hs__nand3_1 _10608_ (.A(net3282),
    .B(net3424),
    .C(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hs__o31ai_1 _10609_ (.A1(_04847_),
    .A2(net3370),
    .A3(net3245),
    .B1(_01985_),
    .Y(_04868_));
 sky130_fd_sc_hs__nor2_2 _10610_ (.A(_04849_),
    .B(net3244),
    .Y(_04869_));
 sky130_fd_sc_hs__nand3b_1 _10611_ (.A_N(_04847_),
    .B(net3200),
    .C(net3684),
    .Y(_04870_));
 sky130_fd_sc_hs__nand2_1 _10612_ (.A(_04868_),
    .B(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hs__inv_2 _10613_ (.A(_04871_),
    .Y(_04872_));
 sky130_fd_sc_hs__buf_1 place2098 (.A(_04591_),
    .X(net2098));
 sky130_fd_sc_hs__nor3_1 _10615_ (.A(_02111_),
    .B(_02108_),
    .C(_04831_),
    .Y(_04874_));
 sky130_fd_sc_hs__inv_1 _10616_ (.A(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hs__nand2_1 _10617_ (.A(_04835_),
    .B(_04822_),
    .Y(_04876_));
 sky130_fd_sc_hs__nor2_4 _10618_ (.A(_04828_),
    .B(net3647),
    .Y(_04877_));
 sky130_fd_sc_hs__nand3_2 _10619_ (.A(net3425),
    .B(net3680),
    .C(_04877_),
    .Y(_04878_));
 sky130_fd_sc_hs__nor3_4 _10620_ (.A(_04875_),
    .B(_04876_),
    .C(_04878_),
    .Y(_04879_));
 sky130_fd_sc_hs__nand3_2 _10621_ (.A(_04819_),
    .B(_04879_),
    .C(_04836_),
    .Y(_04880_));
 sky130_fd_sc_hs__nor3b_4 _10622_ (.A(net3566),
    .B(net3154),
    .C_N(net3429),
    .Y(_04881_));
 sky130_fd_sc_hs__xnor2_2 _10623_ (.A(net3694),
    .B(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hs__xnor2_1 _10624_ (.A(net3695),
    .B(_04869_),
    .Y(_04883_));
 sky130_fd_sc_hs__xnor2_2 _10625_ (.A(_04838_),
    .B(net3697),
    .Y(_04884_));
 sky130_fd_sc_hs__and2_2 _10626_ (.A(_04883_),
    .B(_04884_),
    .X(_04885_));
 sky130_fd_sc_hs__nand2_1 _10627_ (.A(_04848_),
    .B(_04861_),
    .Y(_04886_));
 sky130_fd_sc_hs__nor2_1 _10628_ (.A(_04853_),
    .B(_04859_),
    .Y(_04887_));
 sky130_fd_sc_hs__nor2_1 _10629_ (.A(_04863_),
    .B(_04851_),
    .Y(_04888_));
 sky130_fd_sc_hs__nand2_2 _10630_ (.A(_04887_),
    .B(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hs__nor3_2 _10631_ (.A(net3367),
    .B(_04886_),
    .C(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hs__nor3_1 _10632_ (.A(net3659),
    .B(_02006_),
    .C(_04845_),
    .Y(_04891_));
 sky130_fd_sc_hs__nand2_1 _10633_ (.A(net3198),
    .B(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hs__xnor2_1 _10634_ (.A(net3693),
    .B(_04892_),
    .Y(_04893_));
 sky130_fd_sc_hs__inv_1 _10635_ (.A(_04893_),
    .Y(_04894_));
 sky130_fd_sc_hs__nand3_2 _10636_ (.A(_04885_),
    .B(_04882_),
    .C(_04894_),
    .Y(_04895_));
 sky130_fd_sc_hs__nor2_1 _10637_ (.A(net3638),
    .B(_04878_),
    .Y(_04896_));
 sky130_fd_sc_hs__nand2_1 _10638_ (.A(net3243),
    .B(net3638),
    .Y(_04897_));
 sky130_fd_sc_hs__inv_1 _10639_ (.A(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hs__nor2_1 _10640_ (.A(_04896_),
    .B(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hs__inv_2 _10641_ (.A(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hs__xnor2_4 _10642_ (.A(_04828_),
    .B(net3683),
    .Y(_04901_));
 sky130_fd_sc_hs__nor2_1 _10643_ (.A(net3688),
    .B(_00228_),
    .Y(_04902_));
 sky130_fd_sc_hs__nor2_1 _10644_ (.A(_04902_),
    .B(net5076),
    .Y(_04903_));
 sky130_fd_sc_hs__xnor2_1 _10645_ (.A(_02058_),
    .B(_04857_),
    .Y(_04904_));
 sky130_fd_sc_hs__nor2_1 _10646_ (.A(_04903_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hs__nand2_1 _10647_ (.A(_04905_),
    .B(net3498),
    .Y(_04906_));
 sky130_fd_sc_hs__nor2_1 _10648_ (.A(net3279),
    .B(_04906_),
    .Y(_04907_));
 sky130_fd_sc_hs__xnor2_1 _10649_ (.A(net3570),
    .B(_04858_),
    .Y(_04908_));
 sky130_fd_sc_hs__nand2_1 _10650_ (.A(_04907_),
    .B(net3317),
    .Y(_04909_));
 sky130_fd_sc_hs__inv_1 _10651_ (.A(net3151),
    .Y(_04910_));
 sky130_fd_sc_hs__xnor2_1 _10652_ (.A(net3677),
    .B(net3281),
    .Y(_04911_));
 sky130_fd_sc_hs__xnor2_1 _10653_ (.A(net3680),
    .B(_04859_),
    .Y(_04912_));
 sky130_fd_sc_hs__xnor2_1 _10654_ (.A(net3681),
    .B(_04829_),
    .Y(_04913_));
 sky130_fd_sc_hs__nor2b_2 _10655_ (.A(_04912_),
    .B_N(_04913_),
    .Y(_04914_));
 sky130_fd_sc_hs__nand4_1 _10656_ (.A(net3054),
    .B(_04910_),
    .C(net3241),
    .D(net3197),
    .Y(_04915_));
 sky130_fd_sc_hs__nor2_1 _10657_ (.A(net3366),
    .B(net3243),
    .Y(_04916_));
 sky130_fd_sc_hs__xnor2_1 _10658_ (.A(net3640),
    .B(_04916_),
    .Y(_04917_));
 sky130_fd_sc_hs__xnor2_1 _10659_ (.A(net3709),
    .B(_04889_),
    .Y(_04918_));
 sky130_fd_sc_hs__nor2_1 _10660_ (.A(net3150),
    .B(net3196),
    .Y(_04919_));
 sky130_fd_sc_hs__xnor2_2 _10661_ (.A(net3633),
    .B(_04833_),
    .Y(_04920_));
 sky130_fd_sc_hs__inv_1 _10662_ (.A(net3195),
    .Y(_04921_));
 sky130_fd_sc_hs__xnor2_1 _10663_ (.A(net3636),
    .B(net3282),
    .Y(_04922_));
 sky130_fd_sc_hs__nor2_2 _10664_ (.A(_04921_),
    .B(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hs__nand3b_4 _10665_ (.A_N(_04915_),
    .B(_04919_),
    .C(net3103),
    .Y(_04924_));
 sky130_fd_sc_hs__xnor2_1 _10666_ (.A(net3655),
    .B(net3199),
    .Y(_04925_));
 sky130_fd_sc_hs__o21a_1 _10667_ (.A1(net3368),
    .A2(_04889_),
    .B1(net3658),
    .X(_04926_));
 sky130_fd_sc_hs__nor2_1 _10668_ (.A(net3650),
    .B(_04859_),
    .Y(_04927_));
 sky130_fd_sc_hs__nand4_1 _10669_ (.A(_04927_),
    .B(net3678),
    .C(net3423),
    .D(_04850_),
    .Y(_04928_));
 sky130_fd_sc_hs__nor2_2 _10670_ (.A(net3642),
    .B(_04928_),
    .Y(_04929_));
 sky130_fd_sc_hs__nand2_1 _10671_ (.A(_04929_),
    .B(net3427),
    .Y(_04930_));
 sky130_fd_sc_hs__nor3_1 _10672_ (.A(net3655),
    .B(net3658),
    .C(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hs__nor2_1 _10673_ (.A(_04926_),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hs__nor2_1 _10674_ (.A(_04925_),
    .B(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hs__xnor2_1 _10675_ (.A(net3643),
    .B(_04834_),
    .Y(_04934_));
 sky130_fd_sc_hs__nand2_1 _10676_ (.A(_04929_),
    .B(net3708),
    .Y(_04935_));
 sky130_fd_sc_hs__a22oi_1 _10677_ (.A1(_04929_),
    .A2(net3427),
    .B1(_04935_),
    .B2(net3645),
    .Y(_04936_));
 sky130_fd_sc_hs__nor2_1 _10678_ (.A(net3147),
    .B(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hs__nand3b_4 _10679_ (.A_N(_04924_),
    .B(net3012),
    .C(net3052),
    .Y(_04938_));
 sky130_fd_sc_hs__xnor2_2 _10680_ (.A(_04837_),
    .B(net3704),
    .Y(_04939_));
 sky130_fd_sc_hs__xnor2_1 _10681_ (.A(net3703),
    .B(net3244),
    .Y(_04940_));
 sky130_fd_sc_hs__nor2_2 _10682_ (.A(_04939_),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hs__inv_2 _10683_ (.A(_04941_),
    .Y(_04942_));
 sky130_fd_sc_hs__xnor2_2 _10684_ (.A(net3154),
    .B(net3701),
    .Y(_04943_));
 sky130_fd_sc_hs__xnor2_1 _10685_ (.A(net3699),
    .B(net3198),
    .Y(_04944_));
 sky130_fd_sc_hs__inv_2 _10686_ (.A(_04944_),
    .Y(_04945_));
 sky130_fd_sc_hs__nor2_1 _10687_ (.A(_04943_),
    .B(_04945_),
    .Y(_04946_));
 sky130_fd_sc_hs__inv_1 _10688_ (.A(_04946_),
    .Y(_04947_));
 sky130_fd_sc_hs__nor2_4 _10689_ (.A(_04947_),
    .B(_04942_),
    .Y(_04948_));
 sky130_fd_sc_hs__inv_4 _10690_ (.A(_04948_),
    .Y(_04949_));
 sky130_fd_sc_hs__nor2_1 _10691_ (.A(_04938_),
    .B(net2949),
    .Y(_04950_));
 sky130_fd_sc_hs__nor2_1 _10692_ (.A(net3106),
    .B(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hs__a21oi_1 _10693_ (.A1(net3060),
    .A2(net2975),
    .B1(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hs__xnor2_1 _10694_ (.A(net3015),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hs__inv_1 _10695_ (.A(_04953_),
    .Y(_04954_));
 sky130_fd_sc_hs__nand2_1 _10696_ (.A(_04869_),
    .B(_04846_),
    .Y(_04955_));
 sky130_fd_sc_hs__xnor2_1 _10697_ (.A(net3669),
    .B(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hs__nor2_1 _10698_ (.A(_01965_),
    .B(_01950_),
    .Y(_04957_));
 sky130_fd_sc_hs__and2_1 _10699_ (.A(_04840_),
    .B(_04957_),
    .X(_04958_));
 sky130_fd_sc_hs__nand2_1 _10700_ (.A(_04958_),
    .B(net3429),
    .Y(_04959_));
 sky130_fd_sc_hs__nor2_1 _10701_ (.A(_04959_),
    .B(net3154),
    .Y(_04960_));
 sky130_fd_sc_hs__xnor2_1 _10702_ (.A(net3690),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hs__nand2_1 _10703_ (.A(net3097),
    .B(net3051),
    .Y(_04962_));
 sky130_fd_sc_hs__nand3b_1 _10704_ (.A_N(net3565),
    .B(net3111),
    .C(net3364),
    .Y(_04963_));
 sky130_fd_sc_hs__xnor2_1 _10705_ (.A(net3686),
    .B(_04963_),
    .Y(_04964_));
 sky130_fd_sc_hs__inv_1 _10706_ (.A(_04964_),
    .Y(_04965_));
 sky130_fd_sc_hs__nand3_1 _10707_ (.A(net3422),
    .B(net3693),
    .C(net3690),
    .Y(_04966_));
 sky130_fd_sc_hs__nor2_1 _10708_ (.A(_04966_),
    .B(net3152),
    .Y(_04967_));
 sky130_fd_sc_hs__xnor2_1 _10709_ (.A(net3689),
    .B(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hs__nand3_1 _10710_ (.A(net2973),
    .B(_04872_),
    .C(net3050),
    .Y(_04969_));
 sky130_fd_sc_hs__inv_2 _10711_ (.A(net3056),
    .Y(_04970_));
 sky130_fd_sc_hs__nand2_1 _10712_ (.A(_04911_),
    .B(net3195),
    .Y(_04971_));
 sky130_fd_sc_hs__nor2_1 _10713_ (.A(_00229_),
    .B(net3572),
    .Y(_04972_));
 sky130_fd_sc_hs__inv_2 _10714_ (.A(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hs__nor2_2 _10715_ (.A(_04973_),
    .B(_04903_),
    .Y(_04974_));
 sky130_fd_sc_hs__nor3b_4 _10716_ (.A(_04904_),
    .B(_04901_),
    .C_N(_04974_),
    .Y(_04975_));
 sky130_fd_sc_hs__and2_2 _10717_ (.A(_04975_),
    .B(net3317),
    .X(_04976_));
 sky130_fd_sc_hs__nand3_2 _10718_ (.A(_04900_),
    .B(_04976_),
    .C(_04914_),
    .Y(_04977_));
 sky130_fd_sc_hs__nor2_4 _10719_ (.A(_04977_),
    .B(_04971_),
    .Y(_04978_));
 sky130_fd_sc_hs__nor2_2 _10720_ (.A(_04918_),
    .B(_04934_),
    .Y(_04979_));
 sky130_fd_sc_hs__nor2_1 _10721_ (.A(_04917_),
    .B(_04922_),
    .Y(_04980_));
 sky130_fd_sc_hs__nand3_2 _10722_ (.A(_04978_),
    .B(_04979_),
    .C(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hs__or2_4 _10723_ (.A(net3101),
    .B(_04981_),
    .X(_04982_));
 sky130_fd_sc_hs__inv_1 _10724_ (.A(_04933_),
    .Y(_04983_));
 sky130_fd_sc_hs__nor2_4 _10725_ (.A(_04982_),
    .B(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hs__nor3b_4 _10726_ (.A(_04970_),
    .B(_04949_),
    .C_N(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hs__and2_1 _10727_ (.A(net3057),
    .B(net3153),
    .X(_04986_));
 sky130_fd_sc_hs__and2_2 _10728_ (.A(net3055),
    .B(net3015),
    .X(_04987_));
 sky130_fd_sc_hs__nand3_2 _10729_ (.A(_04985_),
    .B(_04986_),
    .C(_04987_),
    .Y(_04988_));
 sky130_fd_sc_hs__nor3_4 _10730_ (.A(net2855),
    .B(_04969_),
    .C(net3010),
    .Y(_04989_));
 sky130_fd_sc_hs__nand2_1 _10731_ (.A(_04956_),
    .B(_04842_),
    .Y(_04990_));
 sky130_fd_sc_hs__nor3b_1 _10732_ (.A(_04895_),
    .B(_04990_),
    .C_N(_04961_),
    .Y(_04991_));
 sky130_fd_sc_hs__nor3b_4 _10733_ (.A(net3277),
    .B(_04909_),
    .C_N(net3240),
    .Y(_04992_));
 sky130_fd_sc_hs__nand4_2 _10734_ (.A(_04992_),
    .B(_04923_),
    .C(net3241),
    .D(net3054),
    .Y(_04993_));
 sky130_fd_sc_hs__nand3b_4 _10735_ (.A_N(_04993_),
    .B(_04937_),
    .C(net3104),
    .Y(_04994_));
 sky130_fd_sc_hs__nor2_2 _10736_ (.A(net2971),
    .B(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hs__nand4_1 _10737_ (.A(net2947),
    .B(_04991_),
    .C(net2974),
    .D(_04968_),
    .Y(_04996_));
 sky130_fd_sc_hs__nand2_1 _10738_ (.A(_04872_),
    .B(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hs__nand2_2 _10739_ (.A(net2973),
    .B(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hs__nand3_1 _10740_ (.A(net2933),
    .B(net3059),
    .C(net3009),
    .Y(_04999_));
 sky130_fd_sc_hs__nand3_2 _10741_ (.A(_04998_),
    .B(_04989_),
    .C(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hs__nand2_1 _10742_ (.A(_04872_),
    .B(_04988_),
    .Y(_05001_));
 sky130_fd_sc_hs__xnor2_1 _10743_ (.A(net3097),
    .B(_05001_),
    .Y(_05002_));
 sky130_fd_sc_hs__nand2_2 _10744_ (.A(_05000_),
    .B(_05002_),
    .Y(_05003_));
 sky130_fd_sc_hs__inv_2 _10745_ (.A(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hs__o41ai_1 _10746_ (.A1(net2975),
    .A2(net2969),
    .A3(net2949),
    .A4(_04938_),
    .B1(_04872_),
    .Y(_05005_));
 sky130_fd_sc_hs__xnor2_1 _10747_ (.A(net3051),
    .B(net2932),
    .Y(_05006_));
 sky130_fd_sc_hs__nand2_2 _10748_ (.A(_05004_),
    .B(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hs__o21a_1 _10749_ (.A1(net3010),
    .A2(net2855),
    .B1(net3058),
    .X(_05008_));
 sky130_fd_sc_hs__xnor2_2 _10750_ (.A(net3050),
    .B(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hs__nand2_2 _10751_ (.A(net2875),
    .B(_04999_),
    .Y(_05010_));
 sky130_fd_sc_hs__nor2_4 _10752_ (.A(net2840),
    .B(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hs__o211ai_4 _10753_ (.A1(_04954_),
    .A2(_05007_),
    .B1(_05009_),
    .C1(_05011_),
    .Y(_05012_));
 sky130_fd_sc_hs__nand2_1 _10754_ (.A(_04976_),
    .B(net3240),
    .Y(_05013_));
 sky130_fd_sc_hs__nor3_1 _10755_ (.A(net3105),
    .B(net3276),
    .C(net3146),
    .Y(_05014_));
 sky130_fd_sc_hs__nand3_1 _10756_ (.A(net3049),
    .B(net3096),
    .C(net3095),
    .Y(_05015_));
 sky130_fd_sc_hs__nor2_1 _10757_ (.A(net3194),
    .B(net3099),
    .Y(_05016_));
 sky130_fd_sc_hs__inv_2 _10758_ (.A(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hs__clkinv_1 _10759_ (.A(net3053),
    .Y(_05018_));
 sky130_fd_sc_hs__clkinv_1 _10760_ (.A(net3100),
    .Y(_05019_));
 sky130_fd_sc_hs__nor2_1 _10761_ (.A(net3148),
    .B(net3102),
    .Y(_05020_));
 sky130_fd_sc_hs__nand3_1 _10762_ (.A(_05018_),
    .B(_05019_),
    .C(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hs__nor4_2 _10763_ (.A(_04970_),
    .B(net3098),
    .C(_05017_),
    .D(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hs__nand2_1 _10764_ (.A(_04965_),
    .B(_04968_),
    .Y(_05023_));
 sky130_fd_sc_hs__nor2_1 _10765_ (.A(_04962_),
    .B(_05023_),
    .Y(_05024_));
 sky130_fd_sc_hs__nand4_1 _10766_ (.A(_05022_),
    .B(net3005),
    .C(net2970),
    .D(_05024_),
    .Y(_05025_));
 sky130_fd_sc_hs__nor4_2 _10767_ (.A(net3108),
    .B(_05013_),
    .C(net3003),
    .D(_05025_),
    .Y(_05026_));
 sky130_fd_sc_hs__nand2_4 _10768_ (.A(net2874),
    .B(_05010_),
    .Y(_05027_));
 sky130_fd_sc_hs__nand2_2 _10769_ (.A(_05012_),
    .B(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hs__nand2_2 _10770_ (.A(net2856),
    .B(_05028_),
    .Y(_05029_));
 sky130_fd_sc_hs__nand3_2 _10771_ (.A(_05012_),
    .B(net2841),
    .C(_05027_),
    .Y(_05030_));
 sky130_fd_sc_hs__and2_4 _10772_ (.A(_05030_),
    .B(_05029_),
    .X(_05031_));
 sky130_fd_sc_hs__nand2_1 _10773_ (.A(_04985_),
    .B(net3006),
    .Y(_05032_));
 sky130_fd_sc_hs__nand2_1 _10774_ (.A(_05032_),
    .B(net3058),
    .Y(_05033_));
 sky130_fd_sc_hs__xnor2_1 _10775_ (.A(net3055),
    .B(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hs__nand3_2 _10776_ (.A(net2805),
    .B(net2820),
    .C(_05031_),
    .Y(_05035_));
 sky130_fd_sc_hs__inv_1 _10777_ (.A(net2822),
    .Y(_05036_));
 sky130_fd_sc_hs__nand2b_1 _10778_ (.A_N(_05006_),
    .B(net2823),
    .Y(_05037_));
 sky130_fd_sc_hs__nor3_2 _10779_ (.A(_05036_),
    .B(_05037_),
    .C(net2785),
    .Y(_05038_));
 sky130_fd_sc_hs__nand2_2 _10780_ (.A(net2776),
    .B(_05035_),
    .Y(_05039_));
 sky130_fd_sc_hs__nand2_1 _10781_ (.A(net2793),
    .B(net2821),
    .Y(_05040_));
 sky130_fd_sc_hs__nand2_2 _10782_ (.A(net2782),
    .B(_05039_),
    .Y(_05041_));
 sky130_fd_sc_hs__nand2_2 _10783_ (.A(_05041_),
    .B(net2820),
    .Y(_05042_));
 sky130_fd_sc_hs__inv_1 _10784_ (.A(net2820),
    .Y(_05043_));
 sky130_fd_sc_hs__nand3_2 _10785_ (.A(net5060),
    .B(net2812),
    .C(net2783),
    .Y(_05044_));
 sky130_fd_sc_hs__a21oi_1 _10786_ (.A1(net2935),
    .A2(net3014),
    .B1(net3107),
    .Y(_05045_));
 sky130_fd_sc_hs__xnor2_1 _10787_ (.A(net3057),
    .B(_05045_),
    .Y(_05046_));
 sky130_fd_sc_hs__inv_1 _10788_ (.A(_05046_),
    .Y(_05047_));
 sky130_fd_sc_hs__nand3_1 _10789_ (.A(net2736),
    .B(net2741),
    .C(net2854),
    .Y(_05048_));
 sky130_fd_sc_hs__nand2_1 _10790_ (.A(net2777),
    .B(net2784),
    .Y(_05049_));
 sky130_fd_sc_hs__nand2_1 _10791_ (.A(_05042_),
    .B(net2766),
    .Y(_05050_));
 sky130_fd_sc_hs__nand3_1 _10792_ (.A(net2742),
    .B(net2820),
    .C(net2767),
    .Y(_05051_));
 sky130_fd_sc_hs__and2_1 _10793_ (.A(_05050_),
    .B(_05051_),
    .X(_05052_));
 sky130_fd_sc_hs__xnor2_1 _10794_ (.A(_05048_),
    .B(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hs__nand2_1 _10795_ (.A(_05034_),
    .B(_05047_),
    .Y(_05054_));
 sky130_fd_sc_hs__nand2_1 _10796_ (.A(net2805),
    .B(net2841),
    .Y(_05055_));
 sky130_fd_sc_hs__a21oi_1 _10797_ (.A1(_05054_),
    .A2(net2841),
    .B1(net2815),
    .Y(_05056_));
 sky130_fd_sc_hs__o21ai_1 _10798_ (.A1(_05054_),
    .A2(_05055_),
    .B1(_05056_),
    .Y(_05057_));
 sky130_fd_sc_hs__xnor2_1 _10799_ (.A(_05037_),
    .B(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hs__nand2_1 _10800_ (.A(_05058_),
    .B(net2786),
    .Y(_05059_));
 sky130_fd_sc_hs__nand3_1 _10801_ (.A(net2793),
    .B(net2813),
    .C(net2839),
    .Y(_05060_));
 sky130_fd_sc_hs__nand2_1 _10802_ (.A(_05059_),
    .B(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hs__inv_1 _10803_ (.A(_05040_),
    .Y(_05062_));
 sky130_fd_sc_hs__o21ai_1 _10804_ (.A1(_05062_),
    .A2(net2776),
    .B1(_05035_),
    .Y(_05063_));
 sky130_fd_sc_hs__xnor2_2 _10805_ (.A(_05063_),
    .B(_05061_),
    .Y(_05064_));
 sky130_fd_sc_hs__xnor2_2 _10806_ (.A(net2815),
    .B(net5078),
    .Y(_05065_));
 sky130_fd_sc_hs__or2_4 _10807_ (.A(_05065_),
    .B(_05041_),
    .X(_05066_));
 sky130_fd_sc_hs__nor2_2 _10808_ (.A(_05043_),
    .B(_05049_),
    .Y(_05067_));
 sky130_fd_sc_hs__xnor2_1 _10809_ (.A(_05065_),
    .B(_05067_),
    .Y(_05068_));
 sky130_fd_sc_hs__nand2_2 _10810_ (.A(_05041_),
    .B(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hs__nand2_2 _10811_ (.A(_05066_),
    .B(_05069_),
    .Y(_05070_));
 sky130_fd_sc_hs__nor2_2 _10812_ (.A(_05064_),
    .B(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hs__nand4_2 _10813_ (.A(_05042_),
    .B(_05044_),
    .C(net2854),
    .D(net2767),
    .Y(_05072_));
 sky130_fd_sc_hs__nand2_2 _10814_ (.A(_05072_),
    .B(_05071_),
    .Y(_05073_));
 sky130_fd_sc_hs__nand3_1 _10815_ (.A(net2757),
    .B(net2775),
    .C(_05060_),
    .Y(_05074_));
 sky130_fd_sc_hs__o22ai_1 _10816_ (.A1(net2814),
    .A2(net2786),
    .B1(_05040_),
    .B2(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hs__nand2_2 _10817_ (.A(net5065),
    .B(_05075_),
    .Y(_05076_));
 sky130_fd_sc_hs__nand2_2 _10818_ (.A(_05076_),
    .B(_05073_),
    .Y(_05077_));
 sky130_fd_sc_hs__nand2_2 _10819_ (.A(_05053_),
    .B(_05077_),
    .Y(_05078_));
 sky130_fd_sc_hs__nand3_1 _10820_ (.A(_05073_),
    .B(_05076_),
    .C(_05052_),
    .Y(_05079_));
 sky130_fd_sc_hs__nand2_2 _10821_ (.A(_05078_),
    .B(_05079_),
    .Y(_05080_));
 sky130_fd_sc_hs__nand2_1 _10822_ (.A(net2736),
    .B(net2741),
    .Y(_05081_));
 sky130_fd_sc_hs__inv_2 _10823_ (.A(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hs__nand4_1 _10824_ (.A(_05082_),
    .B(net2730),
    .C(net2854),
    .D(net2767),
    .Y(_05083_));
 sky130_fd_sc_hs__nand3_1 _10825_ (.A(net2729),
    .B(net2734),
    .C(net2735),
    .Y(_05084_));
 sky130_fd_sc_hs__nand2_1 _10826_ (.A(_05083_),
    .B(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hs__nand2_2 _10827_ (.A(_05085_),
    .B(_05077_),
    .Y(_05086_));
 sky130_fd_sc_hs__nand3_1 _10828_ (.A(_05073_),
    .B(_05076_),
    .C(net2730),
    .Y(_05087_));
 sky130_fd_sc_hs__nand2_2 _10829_ (.A(_05086_),
    .B(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hs__nor2_4 _10830_ (.A(_05088_),
    .B(_05080_),
    .Y(_05089_));
 sky130_fd_sc_hs__nand2_2 _10831_ (.A(net2854),
    .B(_05077_),
    .Y(_05090_));
 sky130_fd_sc_hs__nand3_1 _10832_ (.A(_05073_),
    .B(net2873),
    .C(_05076_),
    .Y(_05091_));
 sky130_fd_sc_hs__buf_8 place2096 (.A(_05500_),
    .X(net2096));
 sky130_fd_sc_hs__or2_1 _10834_ (.A(net3107),
    .B(_04985_),
    .X(_05093_));
 sky130_fd_sc_hs__xnor2_1 _10835_ (.A(net3153),
    .B(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hs__nand4_2 _10836_ (.A(_05090_),
    .B(_05091_),
    .C(_05094_),
    .D(net2721),
    .Y(_05095_));
 sky130_fd_sc_hs__nand2_2 _10837_ (.A(_05089_),
    .B(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hs__o21ai_1 _10838_ (.A1(net2733),
    .A2(_05084_),
    .B1(net2740),
    .Y(_05097_));
 sky130_fd_sc_hs__nand2_1 _10839_ (.A(_05097_),
    .B(net2710),
    .Y(_05098_));
 sky130_fd_sc_hs__nand2_2 _10840_ (.A(_05096_),
    .B(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hs__xnor2_2 _10841_ (.A(net2692),
    .B(net2722),
    .Y(_05100_));
 sky130_fd_sc_hs__nand3_1 _10842_ (.A(net2693),
    .B(net2701),
    .C(net2837),
    .Y(_05101_));
 sky130_fd_sc_hs__nand2_1 _10843_ (.A(_05101_),
    .B(_05100_),
    .Y(_05102_));
 sky130_fd_sc_hs__nand4_1 _10844_ (.A(net2693),
    .B(net2701),
    .C(net2837),
    .D(net2728),
    .Y(_05103_));
 sky130_fd_sc_hs__nand2_1 _10845_ (.A(_05102_),
    .B(_05103_),
    .Y(_05104_));
 sky130_fd_sc_hs__nand2_2 _10846_ (.A(_05099_),
    .B(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hs__nand3_2 _10847_ (.A(net5089),
    .B(net2700),
    .C(net5064),
    .Y(_05106_));
 sky130_fd_sc_hs__nand2_2 _10848_ (.A(_05106_),
    .B(_05105_),
    .Y(_05107_));
 sky130_fd_sc_hs__inv_1 _10849_ (.A(_05098_),
    .Y(_05108_));
 sky130_fd_sc_hs__o21ai_2 _10850_ (.A1(_05108_),
    .A2(_05089_),
    .B1(net2684),
    .Y(_05109_));
 sky130_fd_sc_hs__nand2_1 _10851_ (.A(net2686),
    .B(_05109_),
    .Y(_05110_));
 sky130_fd_sc_hs__nand2_1 _10852_ (.A(net2693),
    .B(net2701),
    .Y(_05111_));
 sky130_fd_sc_hs__nor2_2 _10853_ (.A(net2728),
    .B(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hs__a21oi_1 _10854_ (.A1(_05112_),
    .A2(net2837),
    .B1(net2686),
    .Y(_05113_));
 sky130_fd_sc_hs__nand2_2 _10855_ (.A(_05099_),
    .B(_05113_),
    .Y(_05114_));
 sky130_fd_sc_hs__nand2_2 _10856_ (.A(_05114_),
    .B(_05110_),
    .Y(_05115_));
 sky130_fd_sc_hs__nor2_2 _10857_ (.A(_05115_),
    .B(_05107_),
    .Y(_05116_));
 sky130_fd_sc_hs__nand3_2 _10858_ (.A(_05096_),
    .B(net2837),
    .C(net2700),
    .Y(_05117_));
 sky130_fd_sc_hs__inv_1 _10859_ (.A(net2837),
    .Y(_05118_));
 sky130_fd_sc_hs__o21ai_1 _10860_ (.A1(_05108_),
    .A2(net2670),
    .B1(_05118_),
    .Y(_05119_));
 sky130_fd_sc_hs__nand2_2 _10861_ (.A(_05119_),
    .B(_05117_),
    .Y(_05120_));
 sky130_fd_sc_hs__xnor2_1 _10862_ (.A(net3008),
    .B(net2903),
    .Y(_05121_));
 sky130_fd_sc_hs__inv_1 _10863_ (.A(net2682),
    .Y(_05122_));
 sky130_fd_sc_hs__nand3_2 _10864_ (.A(_05122_),
    .B(net2871),
    .C(_05120_),
    .Y(_05123_));
 sky130_fd_sc_hs__nand2_2 _10865_ (.A(_05123_),
    .B(_05116_),
    .Y(_05124_));
 sky130_fd_sc_hs__nand3_1 _10866_ (.A(net2683),
    .B(net2694),
    .C(net2702),
    .Y(_05125_));
 sky130_fd_sc_hs__o21ai_2 _10867_ (.A1(_05098_),
    .A2(_05125_),
    .B1(net2685),
    .Y(_05126_));
 sky130_fd_sc_hs__nand2_1 _10868_ (.A(_05126_),
    .B(net2661),
    .Y(_05127_));
 sky130_fd_sc_hs__nand2_2 _10869_ (.A(net2655),
    .B(_05124_),
    .Y(_05128_));
 sky130_fd_sc_hs__nand2_2 _10870_ (.A(net2872),
    .B(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hs__inv_1 _10871_ (.A(net2871),
    .Y(_05130_));
 sky130_fd_sc_hs__o211ai_2 _10872_ (.A1(_05107_),
    .A2(_05115_),
    .B1(_05130_),
    .C1(_05127_),
    .Y(_05131_));
 sky130_fd_sc_hs__a21oi_1 _10873_ (.A1(net2902),
    .A2(net3048),
    .B1(net3108),
    .Y(_05132_));
 sky130_fd_sc_hs__a21oi_1 _10874_ (.A1(net3061),
    .A2(net3002),
    .B1(_05132_),
    .Y(_05133_));
 sky130_fd_sc_hs__xnor2_1 _10875_ (.A(net3098),
    .B(_05133_),
    .Y(_05134_));
 sky130_fd_sc_hs__inv_1 _10876_ (.A(_05134_),
    .Y(_05135_));
 sky130_fd_sc_hs__nand4_2 _10877_ (.A(_05129_),
    .B(_05131_),
    .C(_05135_),
    .D(net2644),
    .Y(_05136_));
 sky130_fd_sc_hs__and2_1 _10878_ (.A(_05126_),
    .B(net2661),
    .X(_05137_));
 sky130_fd_sc_hs__nor2_2 _10879_ (.A(net2638),
    .B(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hs__inv_2 _10880_ (.A(_05107_),
    .Y(_05139_));
 sky130_fd_sc_hs__and2_1 _10881_ (.A(_05123_),
    .B(_05139_),
    .X(_05140_));
 sky130_fd_sc_hs__o21ai_2 _10882_ (.A1(net2653),
    .A2(_05138_),
    .B1(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hs__a21o_1 _10883_ (.A1(_05123_),
    .A2(_05137_),
    .B1(_05139_),
    .X(_05142_));
 sky130_fd_sc_hs__nand2_2 _10884_ (.A(_05142_),
    .B(_05141_),
    .Y(_05143_));
 sky130_fd_sc_hs__xnor2_1 _10885_ (.A(net2837),
    .B(net2682),
    .Y(_05144_));
 sky130_fd_sc_hs__nand2_1 _10886_ (.A(net2656),
    .B(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hs__o21ai_2 _10887_ (.A1(net2682),
    .A2(net2656),
    .B1(_05145_),
    .Y(_05146_));
 sky130_fd_sc_hs__nand2_1 _10888_ (.A(net2644),
    .B(net2871),
    .Y(_05147_));
 sky130_fd_sc_hs__xnor2_1 _10889_ (.A(_05147_),
    .B(_05146_),
    .Y(_05148_));
 sky130_fd_sc_hs__nand2_1 _10890_ (.A(_05128_),
    .B(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hs__nand3_1 _10891_ (.A(_05124_),
    .B(net2637),
    .C(net2655),
    .Y(_05150_));
 sky130_fd_sc_hs__nand2_2 _10892_ (.A(_05149_),
    .B(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hs__nor2_2 _10893_ (.A(_05143_),
    .B(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hs__nand2_2 _10894_ (.A(_05136_),
    .B(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hs__nand2_1 _10895_ (.A(_05123_),
    .B(_05139_),
    .Y(_05154_));
 sky130_fd_sc_hs__o21ai_1 _10896_ (.A1(net2654),
    .A2(_05154_),
    .B1(net2639),
    .Y(_05155_));
 sky130_fd_sc_hs__and2_2 _10897_ (.A(net2617),
    .B(_05155_),
    .X(_05156_));
 sky130_fd_sc_hs__inv_2 _10898_ (.A(net2608),
    .Y(_05157_));
 sky130_fd_sc_hs__nand2_2 _10899_ (.A(_05157_),
    .B(_05153_),
    .Y(_05158_));
 sky130_fd_sc_hs__nand2_2 _10900_ (.A(_05158_),
    .B(net2819),
    .Y(_05159_));
 sky130_fd_sc_hs__nand3_2 _10901_ (.A(_05153_),
    .B(net2836),
    .C(_05157_),
    .Y(_05160_));
 sky130_fd_sc_hs__o21ai_1 _10902_ (.A1(net3011),
    .A2(net2950),
    .B1(net3061),
    .Y(_05161_));
 sky130_fd_sc_hs__xnor2_1 _10903_ (.A(net3099),
    .B(_05161_),
    .Y(_05162_));
 sky130_fd_sc_hs__inv_1 _10904_ (.A(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hs__nand2_2 _10905_ (.A(net2610),
    .B(net2626),
    .Y(_05164_));
 sky130_fd_sc_hs__inv_1 _10906_ (.A(net2600),
    .Y(_05165_));
 sky130_fd_sc_hs__nand4_2 _10907_ (.A(_05159_),
    .B(_05160_),
    .C(_05163_),
    .D(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hs__inv_1 _10908_ (.A(_05151_),
    .Y(_05167_));
 sky130_fd_sc_hs__a21o_1 _10909_ (.A1(_05156_),
    .A2(net2601),
    .B1(_05167_),
    .X(_05168_));
 sky130_fd_sc_hs__and2_1 _10910_ (.A(_05141_),
    .B(_05142_),
    .X(_05169_));
 sky130_fd_sc_hs__o211ai_2 _10911_ (.A1(_05169_),
    .A2(_05156_),
    .B1(_05167_),
    .C1(net2601),
    .Y(_05170_));
 sky130_fd_sc_hs__nand2_2 _10912_ (.A(_05170_),
    .B(_05168_),
    .Y(_05171_));
 sky130_fd_sc_hs__nand2_1 _10913_ (.A(_05129_),
    .B(net2644),
    .Y(_05172_));
 sky130_fd_sc_hs__nand3b_1 _10914_ (.A_N(net2644),
    .B(net5085),
    .C(net2872),
    .Y(_05173_));
 sky130_fd_sc_hs__nand2_1 _10915_ (.A(_05173_),
    .B(_05172_),
    .Y(_05174_));
 sky130_fd_sc_hs__o21ai_1 _10916_ (.A1(net2836),
    .A2(_05164_),
    .B1(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hs__and2_1 _10917_ (.A(_05172_),
    .B(_05173_),
    .X(_05176_));
 sky130_fd_sc_hs__nor2_1 _10918_ (.A(net2836),
    .B(_05164_),
    .Y(_05177_));
 sky130_fd_sc_hs__nand2_1 _10919_ (.A(_05176_),
    .B(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hs__nand2_1 _10920_ (.A(_05175_),
    .B(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hs__nand2_1 _10921_ (.A(_05179_),
    .B(_05158_),
    .Y(_05180_));
 sky130_fd_sc_hs__nand3_1 _10922_ (.A(_05153_),
    .B(net2589),
    .C(_05157_),
    .Y(_05181_));
 sky130_fd_sc_hs__nand2_2 _10923_ (.A(_05181_),
    .B(_05180_),
    .Y(_05182_));
 sky130_fd_sc_hs__nor2_2 _10924_ (.A(_05182_),
    .B(_05171_),
    .Y(_05183_));
 sky130_fd_sc_hs__nand2_2 _10925_ (.A(_05166_),
    .B(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hs__nand2_1 _10926_ (.A(_05170_),
    .B(net2609),
    .Y(_05185_));
 sky130_fd_sc_hs__nand2_1 _10927_ (.A(_05185_),
    .B(net2580),
    .Y(_05186_));
 sky130_fd_sc_hs__nand2_2 _10928_ (.A(_05184_),
    .B(_05186_),
    .Y(_05187_));
 sky130_fd_sc_hs__nand2_2 _10929_ (.A(_05163_),
    .B(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hs__nand3_1 _10930_ (.A(net2536),
    .B(_05162_),
    .C(_05186_),
    .Y(_05189_));
 sky130_fd_sc_hs__xnor2_1 _10931_ (.A(net3194),
    .B(_05132_),
    .Y(_05190_));
 sky130_fd_sc_hs__nand2_1 _10932_ (.A(net2565),
    .B(net2571),
    .Y(_05191_));
 sky130_fd_sc_hs__inv_1 _10933_ (.A(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hs__nand4_2 _10934_ (.A(_05189_),
    .B(_05188_),
    .C(_05190_),
    .D(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hs__xnor2_1 _10935_ (.A(net2819),
    .B(net2600),
    .Y(_05194_));
 sky130_fd_sc_hs__nand2_1 _10936_ (.A(net2572),
    .B(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hs__o21ai_1 _10937_ (.A1(net2600),
    .A2(net2572),
    .B1(_05195_),
    .Y(_05196_));
 sky130_fd_sc_hs__nand3_2 _10938_ (.A(net2565),
    .B(net2571),
    .C(_05163_),
    .Y(_05197_));
 sky130_fd_sc_hs__xnor2_1 _10939_ (.A(_05196_),
    .B(_05197_),
    .Y(_05198_));
 sky130_fd_sc_hs__nand2_1 _10940_ (.A(_05187_),
    .B(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hs__nand3_1 _10941_ (.A(_05184_),
    .B(_05196_),
    .C(_05186_),
    .Y(_05200_));
 sky130_fd_sc_hs__nand2_2 _10942_ (.A(_05199_),
    .B(_05200_),
    .Y(_05201_));
 sky130_fd_sc_hs__nor2_1 _10943_ (.A(net2600),
    .B(_05197_),
    .Y(_05202_));
 sky130_fd_sc_hs__nand2_1 _10944_ (.A(_05202_),
    .B(net2556),
    .Y(_05203_));
 sky130_fd_sc_hs__inv_1 _10945_ (.A(net2555),
    .Y(_05204_));
 sky130_fd_sc_hs__nand2_1 _10946_ (.A(net2557),
    .B(_05204_),
    .Y(_05205_));
 sky130_fd_sc_hs__nand2_1 _10947_ (.A(_05203_),
    .B(_05205_),
    .Y(_05206_));
 sky130_fd_sc_hs__nand2_2 _10948_ (.A(_05206_),
    .B(_05187_),
    .Y(_05207_));
 sky130_fd_sc_hs__nand3_1 _10949_ (.A(net2535),
    .B(net2555),
    .C(_05186_),
    .Y(_05208_));
 sky130_fd_sc_hs__nand2_2 _10950_ (.A(_05207_),
    .B(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hs__nor2_4 _10951_ (.A(_05209_),
    .B(_05201_),
    .Y(_05210_));
 sky130_fd_sc_hs__nand2_2 _10952_ (.A(_05193_),
    .B(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hs__inv_1 _10953_ (.A(net2564),
    .Y(_05212_));
 sky130_fd_sc_hs__nand4_1 _10954_ (.A(_05212_),
    .B(net2557),
    .C(net2546),
    .D(net2570),
    .Y(_05213_));
 sky130_fd_sc_hs__nand3_1 _10955_ (.A(net2534),
    .B(net2578),
    .C(net2579),
    .Y(_05214_));
 sky130_fd_sc_hs__nand2_2 _10956_ (.A(_05213_),
    .B(_05214_),
    .Y(_05215_));
 sky130_fd_sc_hs__inv_1 _10957_ (.A(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hs__nand2_2 _10958_ (.A(_05216_),
    .B(_05211_),
    .Y(_05217_));
 sky130_fd_sc_hs__inv_1 _10959_ (.A(net2515),
    .Y(_05218_));
 sky130_fd_sc_hs__and2_1 _10960_ (.A(net2516),
    .B(_05218_),
    .X(_05219_));
 sky130_fd_sc_hs__nand2_2 _10961_ (.A(_05217_),
    .B(_05219_),
    .Y(_05220_));
 sky130_fd_sc_hs__nand2_1 _10962_ (.A(_05220_),
    .B(net2514),
    .Y(_05221_));
 sky130_fd_sc_hs__nand2_1 _10963_ (.A(_05221_),
    .B(net2492),
    .Y(_05222_));
 sky130_fd_sc_hs__nand3_2 _10964_ (.A(_05216_),
    .B(_05190_),
    .C(_05211_),
    .Y(_05223_));
 sky130_fd_sc_hs__o21bai_1 _10965_ (.A1(net2522),
    .A2(net2504),
    .B1_N(_05190_),
    .Y(_05224_));
 sky130_fd_sc_hs__nand2_2 _10966_ (.A(_05223_),
    .B(_05224_),
    .Y(_05225_));
 sky130_fd_sc_hs__buf_2 place2095 (.A(_05558_),
    .X(net2095));
 sky130_fd_sc_hs__nand2_1 _10968_ (.A(net2950),
    .B(net3061),
    .Y(_05227_));
 sky130_fd_sc_hs__xnor2_1 _10969_ (.A(net3048),
    .B(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hs__nand2_1 _10970_ (.A(net2523),
    .B(net2529),
    .Y(_05229_));
 sky130_fd_sc_hs__inv_1 _10971_ (.A(_05229_),
    .Y(_05230_));
 sky130_fd_sc_hs__nand3_2 _10972_ (.A(_05225_),
    .B(_05228_),
    .C(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hs__xnor2_1 _10973_ (.A(_05163_),
    .B(_05191_),
    .Y(_05232_));
 sky130_fd_sc_hs__nand2_1 _10974_ (.A(net2530),
    .B(_05232_),
    .Y(_05233_));
 sky130_fd_sc_hs__o21ai_2 _10975_ (.A1(net2554),
    .A2(net2530),
    .B1(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hs__nand3_1 _10976_ (.A(net2523),
    .B(net2529),
    .C(_05190_),
    .Y(_05235_));
 sky130_fd_sc_hs__xnor2_1 _10977_ (.A(_05234_),
    .B(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hs__nand2_1 _10978_ (.A(_05217_),
    .B(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hs__nand3_1 _10979_ (.A(net5046),
    .B(_05216_),
    .C(net2513),
    .Y(_05238_));
 sky130_fd_sc_hs__nand2_2 _10980_ (.A(_05238_),
    .B(_05237_),
    .Y(_05239_));
 sky130_fd_sc_hs__inv_1 _10981_ (.A(net2471),
    .Y(_05240_));
 sky130_fd_sc_hs__nand2_1 _10982_ (.A(net2472),
    .B(_05240_),
    .Y(_05241_));
 sky130_fd_sc_hs__o21ai_1 _10983_ (.A1(net2521),
    .A2(net2503),
    .B1(net2516),
    .Y(_05242_));
 sky130_fd_sc_hs__nand2_1 _10984_ (.A(_05242_),
    .B(net2515),
    .Y(_05243_));
 sky130_fd_sc_hs__nand2_2 _10985_ (.A(_05243_),
    .B(_05220_),
    .Y(_05244_));
 sky130_fd_sc_hs__o21ai_1 _10986_ (.A1(net2459),
    .A2(_05241_),
    .B1(net2470),
    .Y(_05245_));
 sky130_fd_sc_hs__nor2_4 _10987_ (.A(_05239_),
    .B(_05244_),
    .Y(_05246_));
 sky130_fd_sc_hs__nand2_2 _10988_ (.A(_05246_),
    .B(_05231_),
    .Y(_05247_));
 sky130_fd_sc_hs__and2_2 _10989_ (.A(_05245_),
    .B(net2449),
    .X(_05248_));
 sky130_fd_sc_hs__nand4_1 _10990_ (.A(net2471),
    .B(net2481),
    .C(_05228_),
    .D(net2502),
    .Y(_05249_));
 sky130_fd_sc_hs__nand2_1 _10991_ (.A(_05249_),
    .B(_05241_),
    .Y(_05250_));
 sky130_fd_sc_hs__nand2_2 _10992_ (.A(_05247_),
    .B(_05222_),
    .Y(_05251_));
 sky130_fd_sc_hs__nand2_2 _10993_ (.A(_05250_),
    .B(_05251_),
    .Y(_05252_));
 sky130_fd_sc_hs__nand3_1 _10994_ (.A(net2448),
    .B(net2459),
    .C(net5103),
    .Y(_05253_));
 sky130_fd_sc_hs__and2_1 _10995_ (.A(_05252_),
    .B(_05253_),
    .X(_05254_));
 sky130_fd_sc_hs__xnor2_1 _10996_ (.A(_05190_),
    .B(_05229_),
    .Y(_05255_));
 sky130_fd_sc_hs__nand2_1 _10997_ (.A(net2488),
    .B(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hs__o21ai_2 _10998_ (.A1(_05229_),
    .A2(net5052),
    .B1(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hs__nand2_1 _10999_ (.A(net2482),
    .B(_05228_),
    .Y(_05258_));
 sky130_fd_sc_hs__xnor2_1 _11000_ (.A(_05258_),
    .B(_05257_),
    .Y(_05259_));
 sky130_fd_sc_hs__nand2_1 _11001_ (.A(_05251_),
    .B(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hs__nand3_1 _11002_ (.A(net5058),
    .B(_05222_),
    .C(net2469),
    .Y(_05261_));
 sky130_fd_sc_hs__nand2_2 _11003_ (.A(_05261_),
    .B(_05260_),
    .Y(_05262_));
 sky130_fd_sc_hs__inv_1 _11004_ (.A(net2427),
    .Y(_05263_));
 sky130_fd_sc_hs__nand2_2 _11005_ (.A(_05251_),
    .B(_05228_),
    .Y(_05264_));
 sky130_fd_sc_hs__inv_1 _11006_ (.A(_05228_),
    .Y(_05265_));
 sky130_fd_sc_hs__nand3_2 _11007_ (.A(net5058),
    .B(_05265_),
    .C(_05222_),
    .Y(_05266_));
 sky130_fd_sc_hs__o21ai_1 _11008_ (.A1(net3148),
    .A2(net2934),
    .B1(net3061),
    .Y(_05267_));
 sky130_fd_sc_hs__xnor2_1 _11009_ (.A(net3001),
    .B(_05267_),
    .Y(_05268_));
 sky130_fd_sc_hs__nand4_2 _11010_ (.A(_05264_),
    .B(_05266_),
    .C(net2870),
    .D(net2483),
    .Y(_05269_));
 sky130_fd_sc_hs__o211ai_1 _11011_ (.A1(_05248_),
    .A2(_05254_),
    .B1(_05263_),
    .C1(net2426),
    .Y(_05270_));
 sky130_fd_sc_hs__nand2_2 _11012_ (.A(_05252_),
    .B(_05253_),
    .Y(_05271_));
 sky130_fd_sc_hs__nand2_1 _11013_ (.A(_05270_),
    .B(net2425),
    .Y(_05272_));
 sky130_fd_sc_hs__nor2_4 _11014_ (.A(_05271_),
    .B(_05262_),
    .Y(_05273_));
 sky130_fd_sc_hs__nand2_2 _11015_ (.A(_05273_),
    .B(_05269_),
    .Y(_05274_));
 sky130_fd_sc_hs__nand2_1 _11016_ (.A(_05272_),
    .B(net2399),
    .Y(_05275_));
 sky130_fd_sc_hs__inv_1 _11017_ (.A(_05248_),
    .Y(_05276_));
 sky130_fd_sc_hs__nand3_2 _11018_ (.A(_05274_),
    .B(net2870),
    .C(_05276_),
    .Y(_05277_));
 sky130_fd_sc_hs__o21bai_1 _11019_ (.A1(_05248_),
    .A2(_05273_),
    .B1_N(net2870),
    .Y(_05278_));
 sky130_fd_sc_hs__nand2_2 _11020_ (.A(_05277_),
    .B(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hs__inv_1 _11021_ (.A(net3148),
    .Y(_05280_));
 sky130_fd_sc_hs__nand2_1 _11022_ (.A(net2968),
    .B(net3061),
    .Y(_05281_));
 sky130_fd_sc_hs__xnor2_1 _11023_ (.A(_05280_),
    .B(_05281_),
    .Y(_05282_));
 sky130_fd_sc_hs__nand2_2 _11024_ (.A(net2433),
    .B(net2440),
    .Y(_05283_));
 sky130_fd_sc_hs__inv_1 _11025_ (.A(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hs__nand3_2 _11026_ (.A(_05279_),
    .B(_05282_),
    .C(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hs__nand2_2 _11027_ (.A(_05274_),
    .B(_05276_),
    .Y(_05286_));
 sky130_fd_sc_hs__inv_1 _11028_ (.A(net2483),
    .Y(_05287_));
 sky130_fd_sc_hs__nand2_1 _11029_ (.A(net2432),
    .B(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hs__nand3_1 _11030_ (.A(net2441),
    .B(_05228_),
    .C(net2483),
    .Y(_05289_));
 sky130_fd_sc_hs__and2_2 _11031_ (.A(_05288_),
    .B(_05289_),
    .X(_05290_));
 sky130_fd_sc_hs__nand3_1 _11032_ (.A(net2432),
    .B(net2440),
    .C(net2870),
    .Y(_05291_));
 sky130_fd_sc_hs__nand2_1 _11033_ (.A(_05290_),
    .B(_05291_),
    .Y(_05292_));
 sky130_fd_sc_hs__nand4_2 _11034_ (.A(net2433),
    .B(net2440),
    .C(net2870),
    .D(_05287_),
    .Y(_05293_));
 sky130_fd_sc_hs__nand2_1 _11035_ (.A(_05293_),
    .B(_05292_),
    .Y(_05294_));
 sky130_fd_sc_hs__nand2_1 _11036_ (.A(_05294_),
    .B(_05286_),
    .Y(_05295_));
 sky130_fd_sc_hs__nand3_1 _11037_ (.A(_05274_),
    .B(net5099),
    .C(_05276_),
    .Y(_05296_));
 sky130_fd_sc_hs__nand2_2 _11038_ (.A(_05296_),
    .B(_05295_),
    .Y(_05297_));
 sky130_fd_sc_hs__inv_1 _11039_ (.A(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hs__nand2_1 _11040_ (.A(_05285_),
    .B(_05298_),
    .Y(_05299_));
 sky130_fd_sc_hs__o21ai_1 _11041_ (.A1(_05248_),
    .A2(net5059),
    .B1(net2426),
    .Y(_05300_));
 sky130_fd_sc_hs__nand2_1 _11042_ (.A(_05300_),
    .B(net2428),
    .Y(_05301_));
 sky130_fd_sc_hs__nand2_2 _11043_ (.A(_05301_),
    .B(_05270_),
    .Y(_05302_));
 sky130_fd_sc_hs__o21ai_1 _11044_ (.A1(_05275_),
    .A2(_05299_),
    .B1(net2382),
    .Y(_05303_));
 sky130_fd_sc_hs__nor2_4 _11045_ (.A(_05302_),
    .B(_05297_),
    .Y(_05304_));
 sky130_fd_sc_hs__nand2_2 _11046_ (.A(_05304_),
    .B(_05285_),
    .Y(_05305_));
 sky130_fd_sc_hs__and2_2 _11047_ (.A(_05303_),
    .B(net2353),
    .X(_05306_));
 sky130_fd_sc_hs__and2_1 _11048_ (.A(_05272_),
    .B(net2399),
    .X(_05307_));
 sky130_fd_sc_hs__inv_1 _11049_ (.A(net2382),
    .Y(_05308_));
 sky130_fd_sc_hs__and2_1 _11050_ (.A(_05285_),
    .B(_05298_),
    .X(_05309_));
 sky130_fd_sc_hs__o21ai_2 _11051_ (.A1(_05307_),
    .A2(_05308_),
    .B1(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hs__a21o_1 _11052_ (.A1(net2373),
    .A2(_05307_),
    .B1(net2358),
    .X(_05311_));
 sky130_fd_sc_hs__nand2_2 _11053_ (.A(_05311_),
    .B(_05310_),
    .Y(_05312_));
 sky130_fd_sc_hs__nand2_2 _11054_ (.A(_05305_),
    .B(_05275_),
    .Y(_05313_));
 sky130_fd_sc_hs__xnor2_1 _11055_ (.A(net2870),
    .B(_05283_),
    .Y(_05314_));
 sky130_fd_sc_hs__nand2_1 _11056_ (.A(net2390),
    .B(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hs__o21ai_1 _11057_ (.A1(net2424),
    .A2(net2390),
    .B1(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hs__nand2_1 _11058_ (.A(net2383),
    .B(_05282_),
    .Y(_05317_));
 sky130_fd_sc_hs__xnor2_1 _11059_ (.A(_05317_),
    .B(_05316_),
    .Y(_05318_));
 sky130_fd_sc_hs__nand2_1 _11060_ (.A(_05313_),
    .B(_05318_),
    .Y(_05319_));
 sky130_fd_sc_hs__nand3_1 _11061_ (.A(net5077),
    .B(net2372),
    .C(_05275_),
    .Y(_05320_));
 sky130_fd_sc_hs__nand2_2 _11062_ (.A(_05320_),
    .B(_05319_),
    .Y(_05321_));
 sky130_fd_sc_hs__nor2_4 _11063_ (.A(_05321_),
    .B(_05312_),
    .Y(_05322_));
 sky130_fd_sc_hs__nand2_2 _11064_ (.A(_05313_),
    .B(_05282_),
    .Y(_05323_));
 sky130_fd_sc_hs__inv_1 _11065_ (.A(_05282_),
    .Y(_05324_));
 sky130_fd_sc_hs__nand3_1 _11066_ (.A(_05305_),
    .B(_05324_),
    .C(_05275_),
    .Y(_05325_));
 sky130_fd_sc_hs__nand2_1 _11067_ (.A(net3061),
    .B(net2948),
    .Y(_05326_));
 sky130_fd_sc_hs__xnor2_1 _11068_ (.A(net3102),
    .B(_05326_),
    .Y(_05327_));
 sky130_fd_sc_hs__inv_1 _11069_ (.A(_05327_),
    .Y(_05328_));
 sky130_fd_sc_hs__nand4_2 _11070_ (.A(_05323_),
    .B(_05325_),
    .C(_05328_),
    .D(net2384),
    .Y(_05329_));
 sky130_fd_sc_hs__o21ai_1 _11071_ (.A1(_05306_),
    .A2(_05322_),
    .B1(net2324),
    .Y(_05330_));
 sky130_fd_sc_hs__nand2_1 _11072_ (.A(_05330_),
    .B(net2325),
    .Y(_05331_));
 sky130_fd_sc_hs__and2_1 _11073_ (.A(_05310_),
    .B(_05311_),
    .X(_05332_));
 sky130_fd_sc_hs__inv_1 _11074_ (.A(net2325),
    .Y(_05333_));
 sky130_fd_sc_hs__o211ai_1 _11075_ (.A1(_05332_),
    .A2(net2337),
    .B1(_05333_),
    .C1(net2324),
    .Y(_05334_));
 sky130_fd_sc_hs__and2_1 _11076_ (.A(_05331_),
    .B(_05334_),
    .X(_05335_));
 sky130_fd_sc_hs__inv_1 _11077_ (.A(_05306_),
    .Y(_05336_));
 sky130_fd_sc_hs__nand2_1 _11078_ (.A(net2324),
    .B(_05333_),
    .Y(_05337_));
 sky130_fd_sc_hs__o21ai_1 _11079_ (.A1(_05336_),
    .A2(_05337_),
    .B1(net2336),
    .Y(_05338_));
 sky130_fd_sc_hs__nand2_2 _11080_ (.A(_05329_),
    .B(_05322_),
    .Y(_05339_));
 sky130_fd_sc_hs__and2_1 _11081_ (.A(_05338_),
    .B(net2308),
    .X(_05340_));
 sky130_fd_sc_hs__nand2_2 _11082_ (.A(_05339_),
    .B(_05336_),
    .Y(_05341_));
 sky130_fd_sc_hs__inv_1 _11083_ (.A(net2384),
    .Y(_05342_));
 sky130_fd_sc_hs__nand2_1 _11084_ (.A(_05323_),
    .B(_05342_),
    .Y(_05343_));
 sky130_fd_sc_hs__nand3_1 _11085_ (.A(net2348),
    .B(_05282_),
    .C(net2384),
    .Y(_05344_));
 sky130_fd_sc_hs__and2_2 _11086_ (.A(_05343_),
    .B(_05344_),
    .X(_05345_));
 sky130_fd_sc_hs__and2_2 _11087_ (.A(net2334),
    .B(net2346),
    .X(_05346_));
 sky130_fd_sc_hs__nand2_1 _11088_ (.A(_05346_),
    .B(_05328_),
    .Y(_05347_));
 sky130_fd_sc_hs__nand2_1 _11089_ (.A(_05347_),
    .B(_05345_),
    .Y(_05348_));
 sky130_fd_sc_hs__nand4_1 _11090_ (.A(net2335),
    .B(net2347),
    .C(_05328_),
    .D(net2371),
    .Y(_05349_));
 sky130_fd_sc_hs__nand2_1 _11091_ (.A(_05348_),
    .B(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hs__nand2_1 _11092_ (.A(_05350_),
    .B(_05341_),
    .Y(_05351_));
 sky130_fd_sc_hs__nand3_1 _11093_ (.A(_05339_),
    .B(_05345_),
    .C(_05336_),
    .Y(_05352_));
 sky130_fd_sc_hs__nand2_2 _11094_ (.A(_05352_),
    .B(_05351_),
    .Y(_05353_));
 sky130_fd_sc_hs__inv_1 _11095_ (.A(net2287),
    .Y(_05354_));
 sky130_fd_sc_hs__nand2_2 _11096_ (.A(_05341_),
    .B(_05328_),
    .Y(_05355_));
 sky130_fd_sc_hs__nand3_2 _11097_ (.A(_05339_),
    .B(_05327_),
    .C(_05336_),
    .Y(_05356_));
 sky130_fd_sc_hs__nand2_1 _11098_ (.A(_04924_),
    .B(net3061),
    .Y(_05357_));
 sky130_fd_sc_hs__xnor2_1 _11099_ (.A(net3147),
    .B(_05357_),
    .Y(_05358_));
 sky130_fd_sc_hs__inv_1 _11100_ (.A(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hs__nand4_2 _11101_ (.A(_05356_),
    .B(_05355_),
    .C(_05359_),
    .D(net2323),
    .Y(_05360_));
 sky130_fd_sc_hs__o211ai_2 _11102_ (.A1(_05335_),
    .A2(_05340_),
    .B1(_05354_),
    .C1(net5051),
    .Y(_05361_));
 sky130_fd_sc_hs__nand2_1 _11103_ (.A(_05331_),
    .B(_05334_),
    .Y(_05362_));
 sky130_fd_sc_hs__nand2_1 _11104_ (.A(net2294),
    .B(_05361_),
    .Y(_05363_));
 sky130_fd_sc_hs__nor2_4 _11105_ (.A(_05362_),
    .B(_05353_),
    .Y(_05364_));
 sky130_fd_sc_hs__nand2_2 _11106_ (.A(_05360_),
    .B(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hs__and2_2 _11107_ (.A(_05363_),
    .B(net2271),
    .X(_05366_));
 sky130_fd_sc_hs__o21ai_1 _11108_ (.A1(_05340_),
    .A2(_05364_),
    .B1(net5051),
    .Y(_05367_));
 sky130_fd_sc_hs__nand2_1 _11109_ (.A(net2288),
    .B(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hs__and2_1 _11110_ (.A(_05368_),
    .B(_05361_),
    .X(_05369_));
 sky130_fd_sc_hs__nand3_1 _11111_ (.A(_05355_),
    .B(_05356_),
    .C(net2323),
    .Y(_05370_));
 sky130_fd_sc_hs__nand2_1 _11112_ (.A(_05364_),
    .B(_05370_),
    .Y(_05371_));
 sky130_fd_sc_hs__inv_1 _11113_ (.A(_05340_),
    .Y(_05372_));
 sky130_fd_sc_hs__nand3_1 _11114_ (.A(_05371_),
    .B(_05359_),
    .C(_05372_),
    .Y(_05373_));
 sky130_fd_sc_hs__o21ai_1 _11115_ (.A1(_05340_),
    .A2(_05364_),
    .B1(_05358_),
    .Y(_05374_));
 sky130_fd_sc_hs__nand2_2 _11116_ (.A(_05374_),
    .B(_05373_),
    .Y(_05375_));
 sky130_fd_sc_hs__inv_1 _11117_ (.A(net2972),
    .Y(_05376_));
 sky130_fd_sc_hs__o31ai_1 _11118_ (.A1(net3150),
    .A2(net3239),
    .A3(_05376_),
    .B1(net3061),
    .Y(_05377_));
 sky130_fd_sc_hs__xnor2_1 _11119_ (.A(net3196),
    .B(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hs__inv_1 _11120_ (.A(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hs__nand2_1 _11121_ (.A(net2296),
    .B(net2302),
    .Y(_05380_));
 sky130_fd_sc_hs__inv_1 _11122_ (.A(net2286),
    .Y(_05381_));
 sky130_fd_sc_hs__nand3_2 _11123_ (.A(_05381_),
    .B(_05379_),
    .C(_05375_),
    .Y(_05382_));
 sky130_fd_sc_hs__xnor2_1 _11124_ (.A(net2323),
    .B(_05355_),
    .Y(_05383_));
 sky130_fd_sc_hs__nand3_1 _11125_ (.A(net2296),
    .B(net2302),
    .C(_05359_),
    .Y(_05384_));
 sky130_fd_sc_hs__nand2_1 _11126_ (.A(_05383_),
    .B(_05384_),
    .Y(_05385_));
 sky130_fd_sc_hs__nand2_1 _11127_ (.A(net2335),
    .B(net2347),
    .Y(_05386_));
 sky130_fd_sc_hs__nand4_1 _11128_ (.A(net2295),
    .B(net2301),
    .C(_05359_),
    .D(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hs__nand2_1 _11129_ (.A(_05385_),
    .B(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hs__nand2_2 _11130_ (.A(_05372_),
    .B(_05365_),
    .Y(_05389_));
 sky130_fd_sc_hs__nand2_2 _11131_ (.A(_05388_),
    .B(_05389_),
    .Y(_05390_));
 sky130_fd_sc_hs__nand3_2 _11132_ (.A(_05365_),
    .B(_05372_),
    .C(_05383_),
    .Y(_05391_));
 sky130_fd_sc_hs__and2_1 _11133_ (.A(_05390_),
    .B(_05391_),
    .X(_05392_));
 sky130_fd_sc_hs__nand2_1 _11134_ (.A(_05382_),
    .B(_05392_),
    .Y(_05393_));
 sky130_fd_sc_hs__o21bai_2 _11135_ (.A1(_05366_),
    .A2(_05369_),
    .B1_N(_05393_),
    .Y(_05394_));
 sky130_fd_sc_hs__nand2_2 _11136_ (.A(_05368_),
    .B(_05361_),
    .Y(_05395_));
 sky130_fd_sc_hs__nand2_1 _11137_ (.A(_05394_),
    .B(net2259),
    .Y(_05396_));
 sky130_fd_sc_hs__nand2_2 _11138_ (.A(_05391_),
    .B(_05390_),
    .Y(_05397_));
 sky130_fd_sc_hs__nor2_4 _11139_ (.A(_05395_),
    .B(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hs__nand2_2 _11140_ (.A(_05398_),
    .B(_05382_),
    .Y(_05399_));
 sky130_fd_sc_hs__nand2_4 _11141_ (.A(_05396_),
    .B(net2233),
    .Y(_05400_));
 sky130_fd_sc_hs__nand2_1 _11142_ (.A(net2260),
    .B(net2275),
    .Y(_05401_));
 sky130_fd_sc_hs__nand3_1 _11143_ (.A(_05392_),
    .B(_05401_),
    .C(_05369_),
    .Y(_05402_));
 sky130_fd_sc_hs__nand2_1 _11144_ (.A(_05363_),
    .B(net2271),
    .Y(_05403_));
 sky130_fd_sc_hs__nand3_1 _11145_ (.A(_05402_),
    .B(_05379_),
    .C(_05403_),
    .Y(_05404_));
 sky130_fd_sc_hs__o21ai_1 _11146_ (.A1(_05366_),
    .A2(_05398_),
    .B1(_05378_),
    .Y(_05405_));
 sky130_fd_sc_hs__nand2_2 _11147_ (.A(_05404_),
    .B(_05405_),
    .Y(_05406_));
 sky130_fd_sc_hs__nand2_1 _11148_ (.A(net3062),
    .B(net3004),
    .Y(_05407_));
 sky130_fd_sc_hs__xnor2_1 _11149_ (.A(net3150),
    .B(_05407_),
    .Y(_05408_));
 sky130_fd_sc_hs__inv_1 _11150_ (.A(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hs__nand3_2 _11151_ (.A(_05406_),
    .B(_05409_),
    .C(net2261),
    .Y(_05410_));
 sky130_fd_sc_hs__nand2_2 _11152_ (.A(_05399_),
    .B(_05403_),
    .Y(_05411_));
 sky130_fd_sc_hs__nand2_1 _11153_ (.A(_05375_),
    .B(_05379_),
    .Y(_05412_));
 sky130_fd_sc_hs__xnor2_1 _11154_ (.A(_05359_),
    .B(_05380_),
    .Y(_05413_));
 sky130_fd_sc_hs__nand2_1 _11155_ (.A(_05389_),
    .B(_05413_),
    .Y(_05414_));
 sky130_fd_sc_hs__o21ai_1 _11156_ (.A1(net2286),
    .A2(_05389_),
    .B1(_05414_),
    .Y(_05415_));
 sky130_fd_sc_hs__xnor2_1 _11157_ (.A(_05412_),
    .B(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hs__nand2_2 _11158_ (.A(_05411_),
    .B(_05416_),
    .Y(_05417_));
 sky130_fd_sc_hs__nand3_1 _11159_ (.A(_05399_),
    .B(_05403_),
    .C(_05415_),
    .Y(_05418_));
 sky130_fd_sc_hs__nand2_2 _11160_ (.A(_05418_),
    .B(_05417_),
    .Y(_05419_));
 sky130_fd_sc_hs__inv_1 _11161_ (.A(net2209),
    .Y(_05420_));
 sky130_fd_sc_hs__nand2_1 _11162_ (.A(net2221),
    .B(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hs__o21ai_2 _11163_ (.A1(_05366_),
    .A2(_05398_),
    .B1(_05382_),
    .Y(_05422_));
 sky130_fd_sc_hs__nand2_1 _11164_ (.A(net2253),
    .B(_05422_),
    .Y(_05423_));
 sky130_fd_sc_hs__nand2_2 _11165_ (.A(_05423_),
    .B(_05394_),
    .Y(_05424_));
 sky130_fd_sc_hs__o21ai_1 _11166_ (.A1(net2222),
    .A2(_05421_),
    .B1(net2220),
    .Y(_05425_));
 sky130_fd_sc_hs__nor2_2 _11167_ (.A(_05424_),
    .B(_05419_),
    .Y(_05426_));
 sky130_fd_sc_hs__nand2_2 _11168_ (.A(_05426_),
    .B(_05410_),
    .Y(_05427_));
 sky130_fd_sc_hs__and2_2 _11169_ (.A(_05425_),
    .B(net5068),
    .X(_05428_));
 sky130_fd_sc_hs__nand4_1 _11170_ (.A(net2209),
    .B(net2229),
    .C(_05409_),
    .D(net2261),
    .Y(_05429_));
 sky130_fd_sc_hs__nand2_1 _11171_ (.A(_05429_),
    .B(_05421_),
    .Y(_05430_));
 sky130_fd_sc_hs__nand2_2 _11172_ (.A(_05427_),
    .B(_05400_),
    .Y(_05431_));
 sky130_fd_sc_hs__nand2_2 _11173_ (.A(net5050),
    .B(_05430_),
    .Y(_05432_));
 sky130_fd_sc_hs__nand3_2 _11174_ (.A(net5068),
    .B(_05400_),
    .C(net2209),
    .Y(_05433_));
 sky130_fd_sc_hs__and2_1 _11175_ (.A(_05432_),
    .B(_05433_),
    .X(_05434_));
 sky130_fd_sc_hs__xnor2_1 _11176_ (.A(_05378_),
    .B(net2261),
    .Y(_05435_));
 sky130_fd_sc_hs__nand2_1 _11177_ (.A(net2228),
    .B(_05435_),
    .Y(_05436_));
 sky130_fd_sc_hs__nand3_1 _11178_ (.A(net2233),
    .B(net2261),
    .C(net2258),
    .Y(_05437_));
 sky130_fd_sc_hs__nand2_1 _11179_ (.A(_05436_),
    .B(_05437_),
    .Y(_05438_));
 sky130_fd_sc_hs__nand2_1 _11180_ (.A(net2229),
    .B(_05409_),
    .Y(_05439_));
 sky130_fd_sc_hs__xnor2_1 _11181_ (.A(_05439_),
    .B(_05438_),
    .Y(_05440_));
 sky130_fd_sc_hs__nand2_1 _11182_ (.A(net5050),
    .B(_05440_),
    .Y(_05441_));
 sky130_fd_sc_hs__nand3_1 _11183_ (.A(_05427_),
    .B(net2208),
    .C(_05400_),
    .Y(_05442_));
 sky130_fd_sc_hs__nand2_2 _11184_ (.A(_05441_),
    .B(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hs__inv_2 _11185_ (.A(net2172),
    .Y(_05444_));
 sky130_fd_sc_hs__nand2_2 _11186_ (.A(_05431_),
    .B(_05409_),
    .Y(_05445_));
 sky130_fd_sc_hs__nand3_2 _11187_ (.A(net5054),
    .B(_05408_),
    .C(_05400_),
    .Y(_05446_));
 sky130_fd_sc_hs__nand2_1 _11188_ (.A(net3062),
    .B(_05376_),
    .Y(_05447_));
 sky130_fd_sc_hs__xnor2_1 _11189_ (.A(net3239),
    .B(_05447_),
    .Y(_05448_));
 sky130_fd_sc_hs__inv_1 _11190_ (.A(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hs__nand4_2 _11191_ (.A(_05446_),
    .B(_05445_),
    .C(_05449_),
    .D(net2230),
    .Y(_05450_));
 sky130_fd_sc_hs__o211ai_2 _11192_ (.A1(_05428_),
    .A2(_05434_),
    .B1(_05444_),
    .C1(net2171),
    .Y(_05451_));
 sky130_fd_sc_hs__a21o_1 _11193_ (.A1(net2171),
    .A2(_05428_),
    .B1(_05444_),
    .X(_05452_));
 sky130_fd_sc_hs__and2_1 _11194_ (.A(_05451_),
    .B(_05452_),
    .X(_05453_));
 sky130_fd_sc_hs__nand2_2 _11195_ (.A(_05433_),
    .B(_05432_),
    .Y(_05454_));
 sky130_fd_sc_hs__nor2_4 _11196_ (.A(_05454_),
    .B(_05443_),
    .Y(_05455_));
 sky130_fd_sc_hs__nand2_2 _11197_ (.A(_05455_),
    .B(_05450_),
    .Y(_05456_));
 sky130_fd_sc_hs__inv_1 _11198_ (.A(net2155),
    .Y(_05457_));
 sky130_fd_sc_hs__a31oi_2 _11199_ (.A1(net2171),
    .A2(_05444_),
    .A3(_05428_),
    .B1(net2173),
    .Y(_05458_));
 sky130_fd_sc_hs__nor2_2 _11200_ (.A(_05457_),
    .B(_05458_),
    .Y(_05459_));
 sky130_fd_sc_hs__inv_1 _11201_ (.A(_05428_),
    .Y(_05460_));
 sky130_fd_sc_hs__nand2_2 _11202_ (.A(_05460_),
    .B(_05456_),
    .Y(_05461_));
 sky130_fd_sc_hs__and2_2 _11203_ (.A(net2181),
    .B(net2191),
    .X(_05462_));
 sky130_fd_sc_hs__nand2_1 _11204_ (.A(_05462_),
    .B(_05449_),
    .Y(_05463_));
 sky130_fd_sc_hs__inv_1 _11205_ (.A(net2230),
    .Y(_05464_));
 sky130_fd_sc_hs__nand2_1 _11206_ (.A(net2181),
    .B(_05464_),
    .Y(_05465_));
 sky130_fd_sc_hs__nand3_1 _11207_ (.A(net2192),
    .B(_05409_),
    .C(net2230),
    .Y(_05466_));
 sky130_fd_sc_hs__and2_2 _11208_ (.A(_05465_),
    .B(_05466_),
    .X(_05467_));
 sky130_fd_sc_hs__nand2_1 _11209_ (.A(_05463_),
    .B(_05467_),
    .Y(_05468_));
 sky130_fd_sc_hs__nand4_1 _11210_ (.A(net2181),
    .B(net5094),
    .C(_05449_),
    .D(net2219),
    .Y(_05469_));
 sky130_fd_sc_hs__nand2_2 _11211_ (.A(_05468_),
    .B(_05469_),
    .Y(_05470_));
 sky130_fd_sc_hs__nand2_2 _11212_ (.A(_05461_),
    .B(_05470_),
    .Y(_05471_));
 sky130_fd_sc_hs__nand3_1 _11213_ (.A(_05456_),
    .B(_05467_),
    .C(_05460_),
    .Y(_05472_));
 sky130_fd_sc_hs__nand2_2 _11214_ (.A(_05472_),
    .B(_05471_),
    .Y(_05473_));
 sky130_fd_sc_hs__inv_2 _11215_ (.A(net2133),
    .Y(_05474_));
 sky130_fd_sc_hs__nand2_2 _11216_ (.A(_05461_),
    .B(_05449_),
    .Y(_05475_));
 sky130_fd_sc_hs__nand3_2 _11217_ (.A(_05456_),
    .B(_05448_),
    .C(_05460_),
    .Y(_05476_));
 sky130_fd_sc_hs__nand2_1 _11218_ (.A(net3062),
    .B(net3013),
    .Y(_05477_));
 sky130_fd_sc_hs__xnor2_1 _11219_ (.A(net3149),
    .B(_05477_),
    .Y(_05478_));
 sky130_fd_sc_hs__inv_1 _11220_ (.A(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hs__nand4_2 _11221_ (.A(_05475_),
    .B(_05476_),
    .C(_05479_),
    .D(net2170),
    .Y(_05480_));
 sky130_fd_sc_hs__o211ai_2 _11222_ (.A1(_05453_),
    .A2(_05459_),
    .B1(_05474_),
    .C1(net5074),
    .Y(_05481_));
 sky130_fd_sc_hs__a21o_1 _11223_ (.A1(_05480_),
    .A2(_05459_),
    .B1(_05474_),
    .X(_05482_));
 sky130_fd_sc_hs__nand2_2 _11224_ (.A(_05482_),
    .B(_05481_),
    .Y(_05483_));
 sky130_fd_sc_hs__nand2_2 _11225_ (.A(_05452_),
    .B(_05451_),
    .Y(_05484_));
 sky130_fd_sc_hs__nor2_4 _11226_ (.A(_05484_),
    .B(_05473_),
    .Y(_05485_));
 sky130_fd_sc_hs__nand2_2 _11227_ (.A(_05480_),
    .B(_05485_),
    .Y(_05486_));
 sky130_fd_sc_hs__or2_4 _11228_ (.A(_05457_),
    .B(_05458_),
    .X(_05487_));
 sky130_fd_sc_hs__nand2_2 _11229_ (.A(_05486_),
    .B(_05487_),
    .Y(_05488_));
 sky130_fd_sc_hs__nand2_1 _11230_ (.A(net2182),
    .B(net5093),
    .Y(_05489_));
 sky130_fd_sc_hs__nand2_1 _11231_ (.A(_05475_),
    .B(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hs__nor2_1 _11232_ (.A(_05448_),
    .B(_05489_),
    .Y(_05491_));
 sky130_fd_sc_hs__nand2_1 _11233_ (.A(net2151),
    .B(_05491_),
    .Y(_05492_));
 sky130_fd_sc_hs__and2_2 _11234_ (.A(_05490_),
    .B(_05492_),
    .X(_05493_));
 sky130_fd_sc_hs__nand3_1 _11235_ (.A(net2143),
    .B(net2149),
    .C(_05479_),
    .Y(_05494_));
 sky130_fd_sc_hs__nand2_1 _11236_ (.A(_05494_),
    .B(_05493_),
    .Y(_05495_));
 sky130_fd_sc_hs__nand4_1 _11237_ (.A(net2143),
    .B(net2149),
    .C(_05479_),
    .D(net2169),
    .Y(_05496_));
 sky130_fd_sc_hs__nand2_1 _11238_ (.A(_05495_),
    .B(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hs__nand2_1 _11239_ (.A(_05497_),
    .B(_05488_),
    .Y(_05498_));
 sky130_fd_sc_hs__nand3_1 _11240_ (.A(_05486_),
    .B(_05487_),
    .C(_05493_),
    .Y(_05499_));
 sky130_fd_sc_hs__nand2_2 _11241_ (.A(_05499_),
    .B(_05498_),
    .Y(_05500_));
 sky130_fd_sc_hs__nor2_4 _11242_ (.A(_05483_),
    .B(_05500_),
    .Y(_05501_));
 sky130_fd_sc_hs__nand3_1 _11243_ (.A(_05475_),
    .B(_05476_),
    .C(net2170),
    .Y(_05502_));
 sky130_fd_sc_hs__nand2_1 _11244_ (.A(_05502_),
    .B(_05485_),
    .Y(_05503_));
 sky130_fd_sc_hs__nand3_2 _11245_ (.A(_05503_),
    .B(_05479_),
    .C(_05487_),
    .Y(_05504_));
 sky130_fd_sc_hs__o21ai_1 _11246_ (.A1(_05459_),
    .A2(_05485_),
    .B1(_05478_),
    .Y(_05505_));
 sky130_fd_sc_hs__nand2_2 _11247_ (.A(_05504_),
    .B(_05505_),
    .Y(_05506_));
 sky130_fd_sc_hs__buf_1 place2094 (.A(net3793),
    .X(net2094));
 sky130_fd_sc_hs__nand2_1 _11249_ (.A(net3062),
    .B(net3007),
    .Y(_05508_));
 sky130_fd_sc_hs__xnor2_1 _11250_ (.A(net3241),
    .B(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hs__nand2_1 _11251_ (.A(net2143),
    .B(net2150),
    .Y(_05510_));
 sky130_fd_sc_hs__inv_2 _11252_ (.A(_05510_),
    .Y(_05511_));
 sky130_fd_sc_hs__nand3_2 _11253_ (.A(_05511_),
    .B(net2946),
    .C(_05506_),
    .Y(_05512_));
 sky130_fd_sc_hs__nand2_2 _11254_ (.A(_05501_),
    .B(_05512_),
    .Y(_05513_));
 sky130_fd_sc_hs__nand2_1 _11255_ (.A(_05481_),
    .B(net2148),
    .Y(_05514_));
 sky130_fd_sc_hs__nand2_4 _11256_ (.A(_05514_),
    .B(net2121),
    .Y(_05515_));
 sky130_fd_sc_hs__nand2_2 _11257_ (.A(_05515_),
    .B(_05513_),
    .Y(_05516_));
 sky130_fd_sc_hs__nand2_2 _11258_ (.A(_05516_),
    .B(net2946),
    .Y(_05517_));
 sky130_fd_sc_hs__inv_1 _11259_ (.A(net2946),
    .Y(_05518_));
 sky130_fd_sc_hs__nand3_1 _11260_ (.A(_05513_),
    .B(_05518_),
    .C(_05515_),
    .Y(_05519_));
 sky130_fd_sc_hs__or2_1 _11261_ (.A(_04992_),
    .B(net3109),
    .X(_05520_));
 sky130_fd_sc_hs__xnor2_1 _11262_ (.A(net3105),
    .B(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hs__inv_1 _11263_ (.A(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hs__nand4_2 _11264_ (.A(_05517_),
    .B(_05519_),
    .C(_05522_),
    .D(net2108),
    .Y(_05523_));
 sky130_fd_sc_hs__nand2_1 _11265_ (.A(net2115),
    .B(_05479_),
    .Y(_05524_));
 sky130_fd_sc_hs__nand2_1 _11266_ (.A(_05524_),
    .B(_05511_),
    .Y(_05525_));
 sky130_fd_sc_hs__nand3_1 _11267_ (.A(net2115),
    .B(_05479_),
    .C(_05510_),
    .Y(_05526_));
 sky130_fd_sc_hs__nand2_1 _11268_ (.A(_05525_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hs__nand2_1 _11269_ (.A(net2107),
    .B(net2946),
    .Y(_05528_));
 sky130_fd_sc_hs__nand2_1 _11270_ (.A(_05527_),
    .B(_05528_),
    .Y(_05529_));
 sky130_fd_sc_hs__inv_1 _11271_ (.A(net2125),
    .Y(_05530_));
 sky130_fd_sc_hs__nand3_1 _11272_ (.A(_05530_),
    .B(net2142),
    .C(_05478_),
    .Y(_05531_));
 sky130_fd_sc_hs__nand4_1 _11273_ (.A(_05524_),
    .B(_05531_),
    .C(net2946),
    .D(net2132),
    .Y(_05532_));
 sky130_fd_sc_hs__nand2_1 _11274_ (.A(_05529_),
    .B(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hs__nand2_1 _11275_ (.A(_05516_),
    .B(_05533_),
    .Y(_05534_));
 sky130_fd_sc_hs__nand3_1 _11276_ (.A(_05513_),
    .B(_05515_),
    .C(_05527_),
    .Y(_05535_));
 sky130_fd_sc_hs__nand2_2 _11277_ (.A(_05534_),
    .B(_05535_),
    .Y(_05536_));
 sky130_fd_sc_hs__nand4_2 _11278_ (.A(net2106),
    .B(net2946),
    .C(net2096),
    .D(net2124),
    .Y(_05537_));
 sky130_fd_sc_hs__inv_1 _11279_ (.A(net2096),
    .Y(_05538_));
 sky130_fd_sc_hs__nand2_1 _11280_ (.A(_05538_),
    .B(net5088),
    .Y(_05539_));
 sky130_fd_sc_hs__nand2_1 _11281_ (.A(_05539_),
    .B(_05537_),
    .Y(_05540_));
 sky130_fd_sc_hs__nand2_1 _11282_ (.A(_05516_),
    .B(_05540_),
    .Y(_05541_));
 sky130_fd_sc_hs__nand3_1 _11283_ (.A(_05513_),
    .B(_05515_),
    .C(net2097),
    .Y(_05542_));
 sky130_fd_sc_hs__nand2_2 _11284_ (.A(_05542_),
    .B(_05541_),
    .Y(_05543_));
 sky130_fd_sc_hs__nor2_4 _11285_ (.A(_05543_),
    .B(_05536_),
    .Y(_05544_));
 sky130_fd_sc_hs__nand2_2 _11286_ (.A(_05544_),
    .B(_05523_),
    .Y(_05545_));
 sky130_fd_sc_hs__o21ai_1 _11287_ (.A1(_05515_),
    .A2(_05539_),
    .B1(net2116),
    .Y(_05546_));
 sky130_fd_sc_hs__nand2_1 _11288_ (.A(_05546_),
    .B(_05513_),
    .Y(_05547_));
 sky130_fd_sc_hs__nand2_2 _11289_ (.A(_05545_),
    .B(_05547_),
    .Y(_05548_));
 sky130_fd_sc_hs__nand2_2 _11290_ (.A(_05522_),
    .B(_05548_),
    .Y(_05549_));
 sky130_fd_sc_hs__nand3_1 _11291_ (.A(_05545_),
    .B(_05521_),
    .C(_05547_),
    .Y(_05550_));
 sky130_fd_sc_hs__nand2_1 _11292_ (.A(net3062),
    .B(net3145),
    .Y(_05551_));
 sky130_fd_sc_hs__xnor2_1 _11293_ (.A(net3278),
    .B(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hs__inv_1 _11294_ (.A(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hs__nand2_1 _11295_ (.A(net2069),
    .B(net2076),
    .Y(_05554_));
 sky130_fd_sc_hs__inv_1 _11296_ (.A(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hs__nand4_1 _11297_ (.A(_05549_),
    .B(_05550_),
    .C(_05553_),
    .D(_05555_),
    .Y(_05556_));
 sky130_fd_sc_hs__nand2_1 _11298_ (.A(_05517_),
    .B(net2108),
    .Y(_05557_));
 sky130_fd_sc_hs__clkinv_1 _11299_ (.A(net2108),
    .Y(_05558_));
 sky130_fd_sc_hs__nand3_1 _11300_ (.A(net2078),
    .B(net2946),
    .C(_05558_),
    .Y(_05559_));
 sky130_fd_sc_hs__nand2_1 _11301_ (.A(_05557_),
    .B(_05559_),
    .Y(_05560_));
 sky130_fd_sc_hs__nand3_1 _11302_ (.A(net5043),
    .B(net2075),
    .C(_05522_),
    .Y(_05561_));
 sky130_fd_sc_hs__nand2_1 _11303_ (.A(_05560_),
    .B(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hs__nand4_1 _11304_ (.A(net2070),
    .B(net2077),
    .C(_05522_),
    .D(net2095),
    .Y(_05563_));
 sky130_fd_sc_hs__nand2_1 _11305_ (.A(_05562_),
    .B(_05563_),
    .Y(_05564_));
 sky130_fd_sc_hs__nand2_1 _11306_ (.A(_05548_),
    .B(_05564_),
    .Y(_05565_));
 sky130_fd_sc_hs__nand3_1 _11307_ (.A(_05545_),
    .B(_05547_),
    .C(_05560_),
    .Y(_05566_));
 sky130_fd_sc_hs__nand2_2 _11308_ (.A(_05565_),
    .B(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hs__nor2_2 _11309_ (.A(net2095),
    .B(_05561_),
    .Y(_05568_));
 sky130_fd_sc_hs__nand2_1 _11310_ (.A(_05568_),
    .B(net2061),
    .Y(_05569_));
 sky130_fd_sc_hs__inv_1 _11311_ (.A(net2061),
    .Y(_05570_));
 sky130_fd_sc_hs__nand2_1 _11312_ (.A(net2062),
    .B(_05570_),
    .Y(_05571_));
 sky130_fd_sc_hs__nand2_1 _11313_ (.A(_05569_),
    .B(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hs__nand2_1 _11314_ (.A(_05572_),
    .B(_05548_),
    .Y(_05573_));
 sky130_fd_sc_hs__nand3_1 _11315_ (.A(_05545_),
    .B(_05547_),
    .C(net2061),
    .Y(_05574_));
 sky130_fd_sc_hs__nand2_1 _11316_ (.A(_05573_),
    .B(_05574_),
    .Y(_05575_));
 sky130_fd_sc_hs__nor2_2 _11317_ (.A(_05567_),
    .B(_05575_),
    .Y(_05576_));
 sky130_fd_sc_hs__nand2_1 _11318_ (.A(_05576_),
    .B(_05556_),
    .Y(_05577_));
 sky130_fd_sc_hs__o21ai_1 _11319_ (.A1(_05547_),
    .A2(_05571_),
    .B1(net2060),
    .Y(_05578_));
 sky130_fd_sc_hs__nand2_1 _11320_ (.A(_05578_),
    .B(net2049),
    .Y(_05579_));
 sky130_fd_sc_hs__nand2_2 _11321_ (.A(_05577_),
    .B(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hs__nand2_2 _11322_ (.A(_05580_),
    .B(_05553_),
    .Y(_05581_));
 sky130_fd_sc_hs__nand3_1 _11323_ (.A(_05577_),
    .B(_05552_),
    .C(_05579_),
    .Y(_05582_));
 sky130_fd_sc_hs__nand2_1 _11324_ (.A(net3062),
    .B(net3151),
    .Y(_05583_));
 sky130_fd_sc_hs__xnor2_1 _11325_ (.A(net3240),
    .B(_05583_),
    .Y(_05584_));
 sky130_fd_sc_hs__and2_4 _11326_ (.A(net2031),
    .B(_05550_),
    .X(_05585_));
 sky130_fd_sc_hs__nand4_2 _11327_ (.A(_05581_),
    .B(_05582_),
    .C(_05584_),
    .D(net2018),
    .Y(_05586_));
 sky130_fd_sc_hs__nand3_1 _11328_ (.A(_05549_),
    .B(_05550_),
    .C(_05555_),
    .Y(_05587_));
 sky130_fd_sc_hs__nor2_1 _11329_ (.A(_05552_),
    .B(_05587_),
    .Y(_05588_));
 sky130_fd_sc_hs__nor2_1 _11330_ (.A(net2020),
    .B(_05588_),
    .Y(_05589_));
 sky130_fd_sc_hs__nand2_1 _11331_ (.A(_05589_),
    .B(_05580_),
    .Y(_05590_));
 sky130_fd_sc_hs__o21ai_1 _11332_ (.A1(_05579_),
    .A2(_05588_),
    .B1(net2020),
    .Y(_05591_));
 sky130_fd_sc_hs__nand2_1 _11333_ (.A(_05590_),
    .B(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hs__nand2_1 _11334_ (.A(net2033),
    .B(net2059),
    .Y(_05593_));
 sky130_fd_sc_hs__nand3_1 _11335_ (.A(net2043),
    .B(_05522_),
    .C(_05555_),
    .Y(_05594_));
 sky130_fd_sc_hs__nand2_1 _11336_ (.A(_05593_),
    .B(_05594_),
    .Y(_05595_));
 sky130_fd_sc_hs__nand3_1 _11337_ (.A(_05595_),
    .B(_05553_),
    .C(_05585_),
    .Y(_05596_));
 sky130_fd_sc_hs__and2_2 _11338_ (.A(_05593_),
    .B(_05594_),
    .X(_05597_));
 sky130_fd_sc_hs__nand2_2 _11339_ (.A(_05585_),
    .B(_05553_),
    .Y(_05598_));
 sky130_fd_sc_hs__nand2_1 _11340_ (.A(_05598_),
    .B(_05597_),
    .Y(_05599_));
 sky130_fd_sc_hs__nand2_1 _11341_ (.A(_05599_),
    .B(_05596_),
    .Y(_05600_));
 sky130_fd_sc_hs__nand2_1 _11342_ (.A(_05600_),
    .B(_05580_),
    .Y(_05601_));
 sky130_fd_sc_hs__nand3_1 _11343_ (.A(net2000),
    .B(_05597_),
    .C(net2029),
    .Y(_05602_));
 sky130_fd_sc_hs__nand2_2 _11344_ (.A(_05602_),
    .B(_05601_),
    .Y(_05603_));
 sky130_fd_sc_hs__nor2_4 _11345_ (.A(_05603_),
    .B(_05592_),
    .Y(_05604_));
 sky130_fd_sc_hs__nand2_2 _11346_ (.A(_05586_),
    .B(_05604_),
    .Y(_05605_));
 sky130_fd_sc_hs__inv_1 _11347_ (.A(net2030),
    .Y(_05606_));
 sky130_fd_sc_hs__nand3_1 _11348_ (.A(_05589_),
    .B(net2019),
    .C(_05606_),
    .Y(_05607_));
 sky130_fd_sc_hs__o21bai_1 _11349_ (.A1(net2020),
    .A2(net2005),
    .B1_N(net2019),
    .Y(_05608_));
 sky130_fd_sc_hs__nand2_1 _11350_ (.A(_05607_),
    .B(_05608_),
    .Y(_05609_));
 sky130_fd_sc_hs__inv_1 _11351_ (.A(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hs__nand2_2 _11352_ (.A(_05605_),
    .B(_05610_),
    .Y(_05611_));
 sky130_fd_sc_hs__nand2_2 _11353_ (.A(_05611_),
    .B(_05584_),
    .Y(_05612_));
 sky130_fd_sc_hs__inv_1 _11354_ (.A(_05584_),
    .Y(_05613_));
 sky130_fd_sc_hs__nand3_2 _11355_ (.A(_05605_),
    .B(_05613_),
    .C(_05610_),
    .Y(_05614_));
 sky130_fd_sc_hs__inv_1 _11356_ (.A(net3318),
    .Y(_05615_));
 sky130_fd_sc_hs__nor2_1 _11357_ (.A(_04975_),
    .B(net3110),
    .Y(_05616_));
 sky130_fd_sc_hs__xnor2_1 _11358_ (.A(_05615_),
    .B(_05616_),
    .Y(_05617_));
 sky130_fd_sc_hs__nand2_1 _11359_ (.A(net1984),
    .B(net1992),
    .Y(_05618_));
 sky130_fd_sc_hs__inv_1 _11360_ (.A(net1974),
    .Y(_05619_));
 sky130_fd_sc_hs__nand4_2 _11361_ (.A(_05612_),
    .B(_05614_),
    .C(net3000),
    .D(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hs__nand2_1 _11362_ (.A(net2032),
    .B(net2042),
    .Y(_05621_));
 sky130_fd_sc_hs__xnor2_1 _11363_ (.A(_05553_),
    .B(_05621_),
    .Y(_05622_));
 sky130_fd_sc_hs__nand2_1 _11364_ (.A(net1993),
    .B(_05622_),
    .Y(_05623_));
 sky130_fd_sc_hs__o21ai_2 _11365_ (.A1(net2016),
    .A2(net1993),
    .B1(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hs__o21ai_1 _11366_ (.A1(_05613_),
    .A2(_05618_),
    .B1(_05624_),
    .Y(_05625_));
 sky130_fd_sc_hs__nand4_1 _11367_ (.A(net1984),
    .B(net1992),
    .C(_05584_),
    .D(net2017),
    .Y(_05626_));
 sky130_fd_sc_hs__nand2_1 _11368_ (.A(_05625_),
    .B(_05626_),
    .Y(_05627_));
 sky130_fd_sc_hs__nand2_1 _11369_ (.A(_05611_),
    .B(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hs__nand3_1 _11370_ (.A(net1961),
    .B(_05610_),
    .C(net1973),
    .Y(_05629_));
 sky130_fd_sc_hs__nand2_1 _11371_ (.A(_05628_),
    .B(_05629_),
    .Y(_05630_));
 sky130_fd_sc_hs__o21ai_1 _11372_ (.A1(_05609_),
    .A2(net1962),
    .B1(net1977),
    .Y(_05631_));
 sky130_fd_sc_hs__nand2_1 _11373_ (.A(_05631_),
    .B(net1975),
    .Y(_05632_));
 sky130_fd_sc_hs__and2_1 _11374_ (.A(_05590_),
    .B(_05591_),
    .X(_05633_));
 sky130_fd_sc_hs__inv_1 _11375_ (.A(net1975),
    .Y(_05634_));
 sky130_fd_sc_hs__o211ai_1 _11376_ (.A1(_05609_),
    .A2(_05633_),
    .B1(_05634_),
    .C1(net1977),
    .Y(_05635_));
 sky130_fd_sc_hs__nand2_1 _11377_ (.A(_05632_),
    .B(_05635_),
    .Y(_05636_));
 sky130_fd_sc_hs__nor2_2 _11378_ (.A(_05630_),
    .B(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hs__nand2_2 _11379_ (.A(_05637_),
    .B(_05620_),
    .Y(_05638_));
 sky130_fd_sc_hs__nand2_1 _11380_ (.A(_05635_),
    .B(net1976),
    .Y(_05639_));
 sky130_fd_sc_hs__nand2_1 _11381_ (.A(_05639_),
    .B(net1960),
    .Y(_05640_));
 sky130_fd_sc_hs__nand2_2 _11382_ (.A(_05638_),
    .B(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hs__and2_4 _11383_ (.A(net1951),
    .B(net1945),
    .X(_05642_));
 sky130_fd_sc_hs__nand2_2 _11384_ (.A(_05642_),
    .B(net3000),
    .Y(_05643_));
 sky130_fd_sc_hs__nor2_1 _11385_ (.A(net1974),
    .B(net1952),
    .Y(_05644_));
 sky130_fd_sc_hs__xnor2_1 _11386_ (.A(_05584_),
    .B(net1974),
    .Y(_05645_));
 sky130_fd_sc_hs__and2_1 _11387_ (.A(_05611_),
    .B(_05645_),
    .X(_05646_));
 sky130_fd_sc_hs__or2_1 _11388_ (.A(_05644_),
    .B(_05646_),
    .X(_05647_));
 sky130_fd_sc_hs__nand2_1 _11389_ (.A(_05647_),
    .B(_05643_),
    .Y(_05648_));
 sky130_fd_sc_hs__nor2_1 _11390_ (.A(_05644_),
    .B(_05646_),
    .Y(_05649_));
 sky130_fd_sc_hs__nand3_2 _11391_ (.A(_05649_),
    .B(_05642_),
    .C(net3000),
    .Y(_05650_));
 sky130_fd_sc_hs__nand2_1 _11392_ (.A(_05650_),
    .B(_05648_),
    .Y(_05651_));
 sky130_fd_sc_hs__nand2_1 _11393_ (.A(_05651_),
    .B(_05641_),
    .Y(_05652_));
 sky130_fd_sc_hs__nand3_1 _11394_ (.A(_05638_),
    .B(_05640_),
    .C(_05647_),
    .Y(_05653_));
 sky130_fd_sc_hs__nand2_2 _11395_ (.A(_05652_),
    .B(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hs__nand3_2 _11396_ (.A(_05638_),
    .B(net3000),
    .C(_05640_),
    .Y(_05655_));
 sky130_fd_sc_hs__and2_2 _11397_ (.A(_05639_),
    .B(net1960),
    .X(_05656_));
 sky130_fd_sc_hs__inv_1 _11398_ (.A(net3000),
    .Y(_05657_));
 sky130_fd_sc_hs__o21ai_1 _11399_ (.A1(_05656_),
    .A2(_05637_),
    .B1(_05657_),
    .Y(_05658_));
 sky130_fd_sc_hs__nand2_2 _11400_ (.A(_05658_),
    .B(_05655_),
    .Y(_05659_));
 sky130_fd_sc_hs__nand2_1 _11401_ (.A(net3062),
    .B(net3242),
    .Y(_05660_));
 sky130_fd_sc_hs__xnor2_1 _11402_ (.A(net3280),
    .B(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hs__inv_1 _11403_ (.A(_05661_),
    .Y(_05662_));
 sky130_fd_sc_hs__nand4_1 _11404_ (.A(net1895),
    .B(net1907),
    .C(_05662_),
    .D(net1933),
    .Y(_05663_));
 sky130_fd_sc_hs__nand3_2 _11405_ (.A(_05659_),
    .B(_05662_),
    .C(net1933),
    .Y(_05664_));
 sky130_fd_sc_hs__inv_1 _11406_ (.A(net1895),
    .Y(_05665_));
 sky130_fd_sc_hs__nand2_1 _11407_ (.A(net1894),
    .B(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hs__nand2_1 _11408_ (.A(_05663_),
    .B(_05666_),
    .Y(_05667_));
 sky130_fd_sc_hs__and2_1 _11409_ (.A(_05632_),
    .B(_05635_),
    .X(_05668_));
 sky130_fd_sc_hs__inv_1 _11410_ (.A(_05630_),
    .Y(_05669_));
 sky130_fd_sc_hs__o211ai_1 _11411_ (.A1(_05668_),
    .A2(_05656_),
    .B1(_05669_),
    .C1(net1934),
    .Y(_05670_));
 sky130_fd_sc_hs__a21o_1 _11412_ (.A1(_05620_),
    .A2(_05656_),
    .B1(_05669_),
    .X(_05671_));
 sky130_fd_sc_hs__nand2_1 _11413_ (.A(_05671_),
    .B(_05670_),
    .Y(_05672_));
 sky130_fd_sc_hs__nor2_4 _11414_ (.A(_05654_),
    .B(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hs__nand2_2 _11415_ (.A(_05664_),
    .B(_05673_),
    .Y(_05674_));
 sky130_fd_sc_hs__nand2_1 _11416_ (.A(_05670_),
    .B(net1944),
    .Y(_05675_));
 sky130_fd_sc_hs__nand2_1 _11417_ (.A(_05675_),
    .B(net1922),
    .Y(_05676_));
 sky130_fd_sc_hs__nand2_2 _11418_ (.A(_05674_),
    .B(_05676_),
    .Y(_05677_));
 sky130_fd_sc_hs__nand2_1 _11419_ (.A(_05667_),
    .B(net5107),
    .Y(_05678_));
 sky130_fd_sc_hs__nand3_1 _11420_ (.A(net1877),
    .B(_05676_),
    .C(net1895),
    .Y(_05679_));
 sky130_fd_sc_hs__nand2_2 _11421_ (.A(_05678_),
    .B(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hs__nand2_1 _11422_ (.A(net1916),
    .B(net3000),
    .Y(_05681_));
 sky130_fd_sc_hs__nand3_1 _11423_ (.A(net1922),
    .B(_05657_),
    .C(net1943),
    .Y(_05682_));
 sky130_fd_sc_hs__nand2_1 _11424_ (.A(_05681_),
    .B(_05682_),
    .Y(_05683_));
 sky130_fd_sc_hs__nand2_1 _11425_ (.A(net1946),
    .B(net1951),
    .Y(_05684_));
 sky130_fd_sc_hs__xnor2_1 _11426_ (.A(net3000),
    .B(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hs__nand2_1 _11427_ (.A(net1916),
    .B(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hs__o21ai_1 _11428_ (.A1(_05684_),
    .A2(net1916),
    .B1(_05686_),
    .Y(_05687_));
 sky130_fd_sc_hs__o21ai_1 _11429_ (.A1(_05661_),
    .A2(_05683_),
    .B1(_05687_),
    .Y(_05688_));
 sky130_fd_sc_hs__nand4_1 _11430_ (.A(_05681_),
    .B(_05682_),
    .C(_05662_),
    .D(net1932),
    .Y(_05689_));
 sky130_fd_sc_hs__nand2_1 _11431_ (.A(_05688_),
    .B(_05689_),
    .Y(_05690_));
 sky130_fd_sc_hs__nand2_1 _11432_ (.A(_05677_),
    .B(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hs__nand3_1 _11433_ (.A(_05674_),
    .B(_05687_),
    .C(net1906),
    .Y(_05692_));
 sky130_fd_sc_hs__nand2_2 _11434_ (.A(_05691_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hs__nand2_2 _11435_ (.A(_05693_),
    .B(_05680_),
    .Y(_05694_));
 sky130_fd_sc_hs__o21ai_2 _11436_ (.A1(net1905),
    .A2(_05666_),
    .B1(net1915),
    .Y(_05695_));
 sky130_fd_sc_hs__nand2_2 _11437_ (.A(_05695_),
    .B(net5055),
    .Y(_05696_));
 sky130_fd_sc_hs__inv_2 _11438_ (.A(_05696_),
    .Y(_05697_));
 sky130_fd_sc_hs__nand2_2 _11439_ (.A(_05677_),
    .B(_05662_),
    .Y(_05698_));
 sky130_fd_sc_hs__nand3_2 _11440_ (.A(_05674_),
    .B(_05661_),
    .C(_05676_),
    .Y(_05699_));
 sky130_fd_sc_hs__and2_4 _11441_ (.A(_05698_),
    .B(_05699_),
    .X(_05700_));
 sky130_fd_sc_hs__nor2_1 _11442_ (.A(net3275),
    .B(net3110),
    .Y(_05701_));
 sky130_fd_sc_hs__xnor2_1 _11443_ (.A(net3365),
    .B(_05701_),
    .Y(_05702_));
 sky130_fd_sc_hs__nor2_1 _11444_ (.A(net3688),
    .B(net3110),
    .Y(_05703_));
 sky130_fd_sc_hs__a21oi_1 _11445_ (.A1(net3110),
    .A2(net3320),
    .B1(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hs__inv_1 _11446_ (.A(_05704_),
    .Y(_05705_));
 sky130_fd_sc_hs__nor3_1 _11447_ (.A(net3428),
    .B(_05705_),
    .C(net1893),
    .Y(_05706_));
 sky130_fd_sc_hs__nand3_2 _11448_ (.A(_05700_),
    .B(_05702_),
    .C(_05706_),
    .Y(_05707_));
 sky130_fd_sc_hs__o31ai_4 _11449_ (.A1(net5084),
    .A2(_05707_),
    .A3(_05694_),
    .B1(net3062),
    .Y(_05708_));
 sky130_fd_sc_hs__buf_1 place2097 (.A(net2096),
    .X(net2097));
 sky130_fd_sc_hs__bufbuf_8 place2093 (.A(_01755_),
    .X(net2093));
 sky130_fd_sc_hs__buf_1 place2092 (.A(_01763_),
    .X(net2092));
 sky130_fd_sc_hs__buf_1 place2091 (.A(_01766_),
    .X(net2091));
 sky130_fd_sc_hs__o21ai_1 _11454_ (.A1(net3778),
    .A2(net3712),
    .B1(net3785),
    .Y(_05713_));
 sky130_fd_sc_hs__a21oi_4 _11455_ (.A1(net5105),
    .A2(net3778),
    .B1(_05713_),
    .Y(_00525_));
 sky130_fd_sc_hs__inv_1 _11456_ (.A(_05680_),
    .Y(_05714_));
 sky130_fd_sc_hs__nor2_2 _11457_ (.A(_05697_),
    .B(_05714_),
    .Y(_05715_));
 sky130_fd_sc_hs__nor2_1 _11458_ (.A(net3363),
    .B(_05705_),
    .Y(_05716_));
 sky130_fd_sc_hs__nand2_1 _11459_ (.A(_05716_),
    .B(_05702_),
    .Y(_05717_));
 sky130_fd_sc_hs__nand2_2 _11460_ (.A(_05698_),
    .B(_05699_),
    .Y(_05718_));
 sky130_fd_sc_hs__nor2_4 _11461_ (.A(_05718_),
    .B(_05717_),
    .Y(_05719_));
 sky130_fd_sc_hs__nand3_2 _11462_ (.A(_05719_),
    .B(net1907),
    .C(_05693_),
    .Y(_05720_));
 sky130_fd_sc_hs__nand2_2 _11463_ (.A(_05720_),
    .B(net3062),
    .Y(_05721_));
 sky130_fd_sc_hs__o211ai_4 _11464_ (.A1(_05715_),
    .A2(net3110),
    .B1(net3778),
    .C1(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hs__buf_1 place2090 (.A(_01775_),
    .X(net2090));
 sky130_fd_sc_hs__a21oi_1 _11466_ (.A1(net3674),
    .A2(net3634),
    .B1(_05774_),
    .Y(_05724_));
 sky130_fd_sc_hs__and2_2 _11467_ (.A(net5044),
    .B(_05724_),
    .X(_00526_));
 sky130_fd_sc_hs__o21ai_1 _11468_ (.A1(net3778),
    .A2(net3710),
    .B1(net3785),
    .Y(_05725_));
 sky130_fd_sc_hs__a21oi_4 _11469_ (.A1(net5105),
    .A2(net3778),
    .B1(_05725_),
    .Y(_00527_));
 sky130_fd_sc_hs__a21oi_1 _11470_ (.A1(net3674),
    .A2(net3641),
    .B1(_05774_),
    .Y(_05726_));
 sky130_fd_sc_hs__and2_2 _11471_ (.A(net5044),
    .B(_05726_),
    .X(_00528_));
 sky130_fd_sc_hs__o21ai_1 _11472_ (.A1(net3778),
    .A2(net3708),
    .B1(net3785),
    .Y(_05727_));
 sky130_fd_sc_hs__a21oi_4 _11473_ (.A1(net5105),
    .A2(net3778),
    .B1(_05727_),
    .Y(_00529_));
 sky130_fd_sc_hs__a21oi_1 _11474_ (.A1(net3674),
    .A2(net3645),
    .B1(_05774_),
    .Y(_05728_));
 sky130_fd_sc_hs__and2_2 _11475_ (.A(net5044),
    .B(_05728_),
    .X(_00530_));
 sky130_fd_sc_hs__o21ai_1 _11476_ (.A1(net3778),
    .A2(net3706),
    .B1(net3785),
    .Y(_05729_));
 sky130_fd_sc_hs__a21oi_4 _11477_ (.A1(net5105),
    .A2(net3778),
    .B1(_05729_),
    .Y(_00531_));
 sky130_fd_sc_hs__a21oi_1 _11478_ (.A1(_00613_),
    .A2(net3656),
    .B1(_05774_),
    .Y(_05730_));
 sky130_fd_sc_hs__and2_2 _11479_ (.A(net1849),
    .B(_05730_),
    .X(_00532_));
 sky130_fd_sc_hs__o21ai_1 _11480_ (.A1(\u_window_buffer.current_state[2] ),
    .A2(net3704),
    .B1(net3785),
    .Y(_05731_));
 sky130_fd_sc_hs__a21oi_4 _11481_ (.A1(net1853),
    .A2(net3778),
    .B1(_05731_),
    .Y(_00533_));
 sky130_fd_sc_hs__a21oi_1 _11482_ (.A1(net3674),
    .A2(net3654),
    .B1(_05774_),
    .Y(_05732_));
 sky130_fd_sc_hs__and2_2 _11483_ (.A(net1849),
    .B(_05732_),
    .X(_00534_));
 sky130_fd_sc_hs__nand2_1 _11484_ (.A(net3674),
    .B(net3702),
    .Y(_05733_));
 sky130_fd_sc_hs__nand2_1 _11485_ (.A(net3778),
    .B(net3497),
    .Y(_05734_));
 sky130_fd_sc_hs__a21oi_1 _11486_ (.A1(_05733_),
    .A2(_05734_),
    .B1(_05774_),
    .Y(_00535_));
 sky130_fd_sc_hs__o21ai_1 _11487_ (.A1(\u_window_buffer.current_state[2] ),
    .A2(net3701),
    .B1(net3784),
    .Y(_05735_));
 sky130_fd_sc_hs__a21oi_4 _11488_ (.A1(net1853),
    .A2(\u_window_buffer.current_state[2] ),
    .B1(_05735_),
    .Y(_00536_));
 sky130_fd_sc_hs__a21oi_1 _11489_ (.A1(_00613_),
    .A2(net3660),
    .B1(_05774_),
    .Y(_05736_));
 sky130_fd_sc_hs__and2_2 _11490_ (.A(net1849),
    .B(_05736_),
    .X(_00537_));
 sky130_fd_sc_hs__o21ai_1 _11491_ (.A1(\u_window_buffer.current_state[2] ),
    .A2(net3698),
    .B1(net3784),
    .Y(_05737_));
 sky130_fd_sc_hs__a21oi_4 _11492_ (.A1(net1853),
    .A2(\u_window_buffer.current_state[2] ),
    .B1(_05737_),
    .Y(_00538_));
 sky130_fd_sc_hs__a21oi_1 _11493_ (.A1(_00613_),
    .A2(_02010_),
    .B1(_05774_),
    .Y(_05738_));
 sky130_fd_sc_hs__and2_2 _11494_ (.A(net1849),
    .B(_05738_),
    .X(_00539_));
 sky130_fd_sc_hs__o21ai_1 _11495_ (.A1(\u_window_buffer.current_state[2] ),
    .A2(net3694),
    .B1(net3784),
    .Y(_05739_));
 sky130_fd_sc_hs__a21oi_4 _11496_ (.A1(net5105),
    .A2(\u_window_buffer.current_state[2] ),
    .B1(_05739_),
    .Y(_00540_));
 sky130_fd_sc_hs__a21oi_1 _11497_ (.A1(_00613_),
    .A2(net3666),
    .B1(_05774_),
    .Y(_05740_));
 sky130_fd_sc_hs__and2_2 _11498_ (.A(net5044),
    .B(_05740_),
    .X(_00541_));
 sky130_fd_sc_hs__o21ai_1 _11499_ (.A1(\u_window_buffer.current_state[2] ),
    .A2(net3692),
    .B1(net3784),
    .Y(_05741_));
 sky130_fd_sc_hs__a21oi_2 _11500_ (.A1(net1853),
    .A2(\u_window_buffer.current_state[2] ),
    .B1(_05741_),
    .Y(_00542_));
 sky130_fd_sc_hs__a21oi_1 _11501_ (.A1(_00613_),
    .A2(net3670),
    .B1(_05774_),
    .Y(_05742_));
 sky130_fd_sc_hs__and2_2 _11502_ (.A(net5044),
    .B(_05742_),
    .X(_00543_));
 sky130_fd_sc_hs__o21ai_1 _11503_ (.A1(\u_window_buffer.current_state[2] ),
    .A2(net3690),
    .B1(net3784),
    .Y(_05743_));
 sky130_fd_sc_hs__a21oi_4 _11504_ (.A1(net1853),
    .A2(\u_window_buffer.current_state[2] ),
    .B1(_05743_),
    .Y(_00544_));
 sky130_fd_sc_hs__a21oi_1 _11505_ (.A1(_00613_),
    .A2(_01994_),
    .B1(_05774_),
    .Y(_05744_));
 sky130_fd_sc_hs__and2_4 _11506_ (.A(net1849),
    .B(_05744_),
    .X(_00545_));
 sky130_fd_sc_hs__nor2_1 _11507_ (.A(net3674),
    .B(net3319),
    .Y(_05745_));
 sky130_fd_sc_hs__a211oi_1 _11508_ (.A1(net3674),
    .A2(net3568),
    .B1(_05774_),
    .C1(_05745_),
    .Y(_00546_));
 sky130_fd_sc_hs__o21ai_1 _11509_ (.A1(\u_window_buffer.current_state[2] ),
    .A2(net3686),
    .B1(net3784),
    .Y(_05746_));
 sky130_fd_sc_hs__a21oi_4 _11510_ (.A1(net1853),
    .A2(\u_window_buffer.current_state[2] ),
    .B1(_05746_),
    .Y(_00547_));
 sky130_fd_sc_hs__a21oi_1 _11511_ (.A1(net3674),
    .A2(net3664),
    .B1(_05774_),
    .Y(_05747_));
 sky130_fd_sc_hs__and2_1 _11512_ (.A(net5044),
    .B(_05747_),
    .X(_00548_));
 sky130_fd_sc_hs__nor2_1 _11513_ (.A(net3110),
    .B(_05716_),
    .Y(_05748_));
 sky130_fd_sc_hs__xor2_1 _11514_ (.A(_05702_),
    .B(_05748_),
    .X(_05749_));
 sky130_fd_sc_hs__o21ai_1 _11515_ (.A1(net3778),
    .A2(\u_window_buffer.write_ptr[3] ),
    .B1(net3785),
    .Y(_05750_));
 sky130_fd_sc_hs__a21oi_1 _11516_ (.A1(_05749_),
    .A2(net3778),
    .B1(_05750_),
    .Y(_00549_));
 sky130_fd_sc_hs__nand2_1 _11517_ (.A(_05702_),
    .B(net3371),
    .Y(_05751_));
 sky130_fd_sc_hs__nand2_1 _11518_ (.A(_05751_),
    .B(net3062),
    .Y(_05752_));
 sky130_fd_sc_hs__xnor2_4 _11519_ (.A(_05752_),
    .B(net1857),
    .Y(_05753_));
 sky130_fd_sc_hs__o21ai_1 _11520_ (.A1(net3778),
    .A2(net3683),
    .B1(net3785),
    .Y(_05754_));
 sky130_fd_sc_hs__a21oi_1 _11521_ (.A1(net3778),
    .A2(_05753_),
    .B1(_05754_),
    .Y(_00550_));
 sky130_fd_sc_hs__xnor2_1 _11522_ (.A(net1907),
    .B(net1863),
    .Y(_05755_));
 sky130_fd_sc_hs__nor2_2 _11523_ (.A(net3110),
    .B(net1854),
    .Y(_05756_));
 sky130_fd_sc_hs__xor2_1 _11524_ (.A(_05755_),
    .B(_05756_),
    .X(_05757_));
 sky130_fd_sc_hs__o21ai_1 _11525_ (.A1(net3778),
    .A2(net3682),
    .B1(net3785),
    .Y(_05758_));
 sky130_fd_sc_hs__a21oi_1 _11526_ (.A1(net1850),
    .A2(net3778),
    .B1(_05758_),
    .Y(_00551_));
 sky130_fd_sc_hs__nand2_1 _11527_ (.A(net1856),
    .B(net3062),
    .Y(_05759_));
 sky130_fd_sc_hs__xnor2_2 _11528_ (.A(net1859),
    .B(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hs__o21ai_1 _11529_ (.A1(net3778),
    .A2(net3681),
    .B1(net3785),
    .Y(_05761_));
 sky130_fd_sc_hs__a21oi_1 _11530_ (.A1(_05760_),
    .A2(net3778),
    .B1(_05761_),
    .Y(_00552_));
 sky130_fd_sc_hs__nand2_1 _11531_ (.A(net1855),
    .B(net5071),
    .Y(_05762_));
 sky130_fd_sc_hs__nand3_1 _11532_ (.A(net1852),
    .B(net3062),
    .C(net1860),
    .Y(_05763_));
 sky130_fd_sc_hs__o21ai_1 _11533_ (.A1(net3778),
    .A2(net3680),
    .B1(net3785),
    .Y(_05764_));
 sky130_fd_sc_hs__a31oi_2 _11534_ (.A1(_05763_),
    .A2(_05762_),
    .A3(net3778),
    .B1(_05764_),
    .Y(_00553_));
 sky130_fd_sc_hs__nand3_1 _11535_ (.A(net1862),
    .B(net1870),
    .C(net1907),
    .Y(_05765_));
 sky130_fd_sc_hs__o21ai_2 _11536_ (.A1(_05765_),
    .A2(_05694_),
    .B1(net3062),
    .Y(_05766_));
 sky130_fd_sc_hs__nand2_1 _11537_ (.A(_05766_),
    .B(_05752_),
    .Y(_05767_));
 sky130_fd_sc_hs__nand2_1 _11538_ (.A(_05767_),
    .B(net1864),
    .Y(_05768_));
 sky130_fd_sc_hs__nand3_1 _11539_ (.A(_05766_),
    .B(net1858),
    .C(_05752_),
    .Y(_05769_));
 sky130_fd_sc_hs__nand3_2 _11540_ (.A(_05768_),
    .B(_05769_),
    .C(net3778),
    .Y(_05770_));
 sky130_fd_sc_hs__a21oi_1 _11541_ (.A1(net3674),
    .A2(net3638),
    .B1(_05774_),
    .Y(_05771_));
 sky130_fd_sc_hs__and2_2 _11542_ (.A(_05770_),
    .B(_05771_),
    .X(_00554_));
 sky130_fd_sc_hs__a21oi_1 _11543_ (.A1(net3674),
    .A2(net3637),
    .B1(_05774_),
    .Y(_05772_));
 sky130_fd_sc_hs__and2_1 _11544_ (.A(net1849),
    .B(_05772_),
    .X(_00555_));
 sky130_fd_sc_hs__fa_1 _11545_ (.A(\u_fft.sched[31] ),
    .B(\u_fft.sched[56] ),
    .CIN(_00026_),
    .COUT(_00027_),
    .SUM(_00028_));
 sky130_fd_sc_hs__ha_1 _11546_ (.A(\u_fft.sched[54] ),
    .B(_00029_),
    .COUT(_00030_),
    .SUM(_00031_));
 sky130_fd_sc_hs__ha_1 _11547_ (.A(\u_fft.sched[53] ),
    .B(_00032_),
    .COUT(_00033_),
    .SUM(_00034_));
 sky130_fd_sc_hs__ha_1 _11548_ (.A(\u_fft.sched[52] ),
    .B(_00035_),
    .COUT(_00036_),
    .SUM(_00037_));
 sky130_fd_sc_hs__ha_1 _11549_ (.A(\u_fft.sched[51] ),
    .B(_00038_),
    .COUT(_00039_),
    .SUM(_00040_));
 sky130_fd_sc_hs__ha_1 _11550_ (.A(\u_fft.sched[50] ),
    .B(_00041_),
    .COUT(_00042_),
    .SUM(_00043_));
 sky130_fd_sc_hs__ha_1 _11551_ (.A(\u_fft.sched[49] ),
    .B(_00044_),
    .COUT(_00045_),
    .SUM(_00046_));
 sky130_fd_sc_hs__ha_1 _11552_ (.A(\u_fft.sched[48] ),
    .B(_00047_),
    .COUT(_00048_),
    .SUM(_00049_));
 sky130_fd_sc_hs__ha_1 _11553_ (.A(\u_fft.sched[47] ),
    .B(_00050_),
    .COUT(_00051_),
    .SUM(_00052_));
 sky130_fd_sc_hs__ha_1 _11554_ (.A(_00053_),
    .B(_00054_),
    .COUT(_00055_),
    .SUM(_05851_));
 sky130_fd_sc_hs__ha_1 _11555_ (.A(\u_fft.sched[46] ),
    .B(_05851_),
    .COUT(_00056_),
    .SUM(_00057_));
 sky130_fd_sc_hs__ha_1 _11556_ (.A(\u_fft.sched[64] ),
    .B(_00058_),
    .COUT(_00059_),
    .SUM(_00060_));
 sky130_fd_sc_hs__ha_1 _11557_ (.A(\u_fft.sched[63] ),
    .B(_00061_),
    .COUT(_00062_),
    .SUM(_00063_));
 sky130_fd_sc_hs__ha_1 _11558_ (.A(\u_fft.sched[62] ),
    .B(_00064_),
    .COUT(_00065_),
    .SUM(_00066_));
 sky130_fd_sc_hs__ha_1 _11559_ (.A(\u_fft.sched[61] ),
    .B(_00067_),
    .COUT(_00068_),
    .SUM(_00069_));
 sky130_fd_sc_hs__ha_1 _11560_ (.A(\u_fft.sched[60] ),
    .B(_00070_),
    .COUT(_00071_),
    .SUM(_00072_));
 sky130_fd_sc_hs__ha_1 _11561_ (.A(\u_fft.sched[59] ),
    .B(_00073_),
    .COUT(_00074_),
    .SUM(_00075_));
 sky130_fd_sc_hs__ha_1 _11562_ (.A(\u_fft.sched[58] ),
    .B(_00076_),
    .COUT(_00077_),
    .SUM(_00078_));
 sky130_fd_sc_hs__ha_1 _11563_ (.A(\u_fft.sched[57] ),
    .B(_00079_),
    .COUT(_00080_),
    .SUM(_00081_));
 sky130_fd_sc_hs__ha_1 _11564_ (.A(_00082_),
    .B(_00083_),
    .COUT(_00084_),
    .SUM(_00085_));
 sky130_fd_sc_hs__ha_1 _11565_ (.A(\u_fft.sched[56] ),
    .B(_00086_),
    .COUT(_00087_),
    .SUM(_00088_));
 sky130_fd_sc_hs__ha_1 _11566_ (.A(\u_window_buffer.read_ptr[30] ),
    .B(\u_window_buffer.internal_read_ptr[30] ),
    .COUT(_00089_),
    .SUM(_00090_));
 sky130_fd_sc_hs__ha_1 _11567_ (.A(\u_window_buffer.read_ptr[29] ),
    .B(\u_window_buffer.internal_read_ptr[29] ),
    .COUT(_00091_),
    .SUM(_00092_));
 sky130_fd_sc_hs__ha_1 _11568_ (.A(\u_window_buffer.read_ptr[28] ),
    .B(\u_window_buffer.internal_read_ptr[28] ),
    .COUT(_00093_),
    .SUM(_00094_));
 sky130_fd_sc_hs__ha_1 _11569_ (.A(\u_window_buffer.read_ptr[27] ),
    .B(\u_window_buffer.internal_read_ptr[27] ),
    .COUT(_00095_),
    .SUM(_00096_));
 sky130_fd_sc_hs__ha_1 _11570_ (.A(\u_window_buffer.read_ptr[26] ),
    .B(\u_window_buffer.internal_read_ptr[26] ),
    .COUT(_00097_),
    .SUM(_00098_));
 sky130_fd_sc_hs__ha_1 _11571_ (.A(\u_window_buffer.internal_read_ptr[25] ),
    .B(\u_window_buffer.read_ptr[25] ),
    .COUT(_00099_),
    .SUM(_00100_));
 sky130_fd_sc_hs__ha_1 _11572_ (.A(\u_window_buffer.read_ptr[24] ),
    .B(\u_window_buffer.internal_read_ptr[24] ),
    .COUT(_00101_),
    .SUM(_00102_));
 sky130_fd_sc_hs__ha_1 _11573_ (.A(\u_window_buffer.read_ptr[23] ),
    .B(\u_window_buffer.internal_read_ptr[23] ),
    .COUT(_00103_),
    .SUM(_00104_));
 sky130_fd_sc_hs__ha_1 _11574_ (.A(\u_window_buffer.read_ptr[22] ),
    .B(\u_window_buffer.internal_read_ptr[22] ),
    .COUT(_00105_),
    .SUM(_00106_));
 sky130_fd_sc_hs__ha_1 _11575_ (.A(\u_window_buffer.internal_read_ptr[21] ),
    .B(\u_window_buffer.read_ptr[21] ),
    .COUT(_00107_),
    .SUM(_00108_));
 sky130_fd_sc_hs__ha_4 _11576_ (.A(\u_window_buffer.read_ptr[20] ),
    .B(\u_window_buffer.internal_read_ptr[20] ),
    .COUT(_00109_),
    .SUM(_00110_));
 sky130_fd_sc_hs__ha_1 _11577_ (.A(\u_window_buffer.internal_read_ptr[19] ),
    .B(\u_window_buffer.read_ptr[19] ),
    .COUT(_00111_),
    .SUM(_00112_));
 sky130_fd_sc_hs__ha_1 _11578_ (.A(\u_window_buffer.read_ptr[18] ),
    .B(\u_window_buffer.internal_read_ptr[18] ),
    .COUT(_00113_),
    .SUM(_00114_));
 sky130_fd_sc_hs__ha_1 _11579_ (.A(\u_window_buffer.internal_read_ptr[17] ),
    .B(\u_window_buffer.read_ptr[17] ),
    .COUT(_00115_),
    .SUM(_00116_));
 sky130_fd_sc_hs__ha_1 _11580_ (.A(\u_window_buffer.read_ptr[16] ),
    .B(\u_window_buffer.internal_read_ptr[16] ),
    .COUT(_00117_),
    .SUM(_00118_));
 sky130_fd_sc_hs__ha_1 _11581_ (.A(\u_window_buffer.internal_read_ptr[15] ),
    .B(\u_window_buffer.read_ptr[15] ),
    .COUT(_00119_),
    .SUM(_00120_));
 sky130_fd_sc_hs__ha_1 _11582_ (.A(\u_window_buffer.read_ptr[14] ),
    .B(\u_window_buffer.internal_read_ptr[14] ),
    .COUT(_00121_),
    .SUM(_00122_));
 sky130_fd_sc_hs__ha_4 _11583_ (.A(\u_window_buffer.read_ptr[13] ),
    .B(net3772),
    .COUT(_00123_),
    .SUM(_00124_));
 sky130_fd_sc_hs__ha_4 _11584_ (.A(\u_window_buffer.read_ptr[12] ),
    .B(\u_window_buffer.internal_read_ptr[12] ),
    .COUT(_00125_),
    .SUM(_00126_));
 sky130_fd_sc_hs__ha_2 _11585_ (.A(\u_window_buffer.internal_read_ptr[11] ),
    .B(\u_window_buffer.read_ptr[11] ),
    .COUT(_00127_),
    .SUM(_00128_));
 sky130_fd_sc_hs__ha_4 _11586_ (.A(\u_window_buffer.internal_read_ptr[10] ),
    .B(\u_window_buffer.read_ptr[10] ),
    .COUT(_00129_),
    .SUM(_00130_));
 sky130_fd_sc_hs__ha_4 _11587_ (.A(\u_window_buffer.read_ptr[9] ),
    .B(\u_window_buffer.internal_read_ptr[9] ),
    .COUT(_00131_),
    .SUM(_00132_));
 sky130_fd_sc_hs__ha_4 _11588_ (.A(\u_window_buffer.read_ptr[8] ),
    .B(\u_window_buffer.internal_read_ptr[8] ),
    .COUT(_00133_),
    .SUM(_00134_));
 sky130_fd_sc_hs__ha_2 _11589_ (.A(\u_window_buffer.internal_read_ptr[7] ),
    .B(\u_window_buffer.read_ptr[7] ),
    .COUT(_00135_),
    .SUM(_00136_));
 sky130_fd_sc_hs__ha_4 _11590_ (.A(\u_window_buffer.internal_read_ptr[6] ),
    .B(\u_window_buffer.read_ptr[6] ),
    .COUT(_00137_),
    .SUM(_00138_));
 sky130_fd_sc_hs__ha_4 _11591_ (.A(\u_window_buffer.read_ptr[5] ),
    .B(\u_window_buffer.internal_read_ptr[5] ),
    .COUT(_00139_),
    .SUM(_00140_));
 sky130_fd_sc_hs__ha_4 _11592_ (.A(\u_window_buffer.internal_read_ptr[4] ),
    .B(\u_window_buffer.read_ptr[4] ),
    .COUT(_00141_),
    .SUM(_00142_));
 sky130_fd_sc_hs__ha_4 _11593_ (.A(\u_window_buffer.internal_read_ptr[3] ),
    .B(\u_window_buffer.read_ptr[3] ),
    .COUT(_00143_),
    .SUM(_00144_));
 sky130_fd_sc_hs__ha_4 _11594_ (.A(\u_window_buffer.read_ptr[2] ),
    .B(\u_window_buffer.internal_read_ptr[2] ),
    .COUT(_00145_),
    .SUM(_00146_));
 sky130_fd_sc_hs__ha_1 _11595_ (.A(\u_window_buffer.read_ptr[1] ),
    .B(\u_window_buffer.internal_read_ptr[1] ),
    .COUT(_00147_),
    .SUM(_00148_));
 sky130_fd_sc_hs__ha_1 _11596_ (.A(\u_window_buffer.read_ptr[1] ),
    .B(\u_window_buffer.internal_read_ptr[1] ),
    .COUT(_00149_),
    .SUM(_05852_));
 sky130_fd_sc_hs__ha_1 _11597_ (.A(_00150_),
    .B(_00151_),
    .COUT(_00152_),
    .SUM(_00153_));
 sky130_fd_sc_hs__ha_1 _11598_ (.A(net3672),
    .B(_00154_),
    .COUT(_00155_),
    .SUM(_00156_));
 sky130_fd_sc_hs__ha_1 _11599_ (.A(\tx_fifo.write_ptr[0] ),
    .B(\tx_fifo.write_ptr[1] ),
    .COUT(_00157_),
    .SUM(_00158_));
 sky130_fd_sc_hs__ha_1 _11600_ (.A(_00159_),
    .B(_00160_),
    .COUT(_00161_),
    .SUM(_00162_));
 sky130_fd_sc_hs__ha_1 _11601_ (.A(\u_dct.k_ptr[0] ),
    .B(\u_dct.k_ptr[1] ),
    .COUT(_00163_),
    .SUM(_05853_));
 sky130_fd_sc_hs__ha_1 _11602_ (.A(_00164_),
    .B(_00165_),
    .COUT(_00166_),
    .SUM(_00167_));
 sky130_fd_sc_hs__ha_1 _11603_ (.A(\u_dct.n_ptr[0] ),
    .B(\u_dct.n_ptr[1] ),
    .COUT(_00168_),
    .SUM(_05854_));
 sky130_fd_sc_hs__ha_1 _11604_ (.A(_00169_),
    .B(_00170_),
    .COUT(_00171_),
    .SUM(_00172_));
 sky130_fd_sc_hs__ha_1 _11605_ (.A(_00169_),
    .B(\u_fft.sched[41] ),
    .COUT(_00173_),
    .SUM(_05855_));
 sky130_fd_sc_hs__ha_1 _11606_ (.A(\u_fft.sched[40] ),
    .B(_00170_),
    .COUT(_00174_),
    .SUM(_05856_));
 sky130_fd_sc_hs__ha_1 _11607_ (.A(\u_fft.sched[40] ),
    .B(\u_fft.sched[41] ),
    .COUT(_00175_),
    .SUM(_05857_));
 sky130_fd_sc_hs__ha_1 _11608_ (.A(_00176_),
    .B(_00175_),
    .COUT(_00177_),
    .SUM(_00178_));
 sky130_fd_sc_hs__ha_1 _11609_ (.A(\u_fft.sched[42] ),
    .B(_00175_),
    .COUT(_00179_),
    .SUM(_05858_));
 sky130_fd_sc_hs__ha_1 _11610_ (.A(\u_fft.sched[45] ),
    .B(\u_fft.sched[46] ),
    .COUT(_00180_),
    .SUM(_00181_));
 sky130_fd_sc_hs__ha_1 _11611_ (.A(\u_fft.sched[30] ),
    .B(_00182_),
    .COUT(_00183_),
    .SUM(_00184_));
 sky130_fd_sc_hs__ha_1 _11612_ (.A(\u_fft.sched[30] ),
    .B(\u_fft.sched[55] ),
    .COUT(_00026_),
    .SUM(_05859_));
 sky130_fd_sc_hs__ha_1 _11613_ (.A(\u_fft.sched[31] ),
    .B(\u_fft.sched[56] ),
    .COUT(_00185_),
    .SUM(_00186_));
 sky130_fd_sc_hs__ha_1 _11614_ (.A(\u_fft.sched[32] ),
    .B(\u_fft.sched[57] ),
    .COUT(_00187_),
    .SUM(_00188_));
 sky130_fd_sc_hs__ha_1 _11615_ (.A(\u_fft.sched[33] ),
    .B(\u_fft.sched[58] ),
    .COUT(_00189_),
    .SUM(_00190_));
 sky130_fd_sc_hs__ha_1 _11616_ (.A(\u_fft.sched[34] ),
    .B(\u_fft.sched[59] ),
    .COUT(_00191_),
    .SUM(_00192_));
 sky130_fd_sc_hs__ha_1 _11617_ (.A(\u_fft.sched[35] ),
    .B(\u_fft.sched[60] ),
    .COUT(_00193_),
    .SUM(_00194_));
 sky130_fd_sc_hs__ha_1 _11618_ (.A(\u_fft.sched[36] ),
    .B(\u_fft.sched[61] ),
    .COUT(_00195_),
    .SUM(_00196_));
 sky130_fd_sc_hs__ha_1 _11619_ (.A(\u_fft.sched[37] ),
    .B(\u_fft.sched[62] ),
    .COUT(_00197_),
    .SUM(_00198_));
 sky130_fd_sc_hs__ha_1 _11620_ (.A(\u_fft.sched[38] ),
    .B(\u_fft.sched[63] ),
    .COUT(_00199_),
    .SUM(_00200_));
 sky130_fd_sc_hs__ha_1 _11621_ (.A(\u_fft.power_ptr[0] ),
    .B(\u_fft.power_ptr[1] ),
    .COUT(_00201_),
    .SUM(_00202_));
 sky130_fd_sc_hs__ha_1 _11622_ (.A(\u_hamming_window.frame_ptr[0] ),
    .B(\u_hamming_window.frame_ptr[1] ),
    .COUT(_00203_),
    .SUM(_00204_));
 sky130_fd_sc_hs__ha_1 _11623_ (.A(_00205_),
    .B(_00206_),
    .COUT(_00207_),
    .SUM(_00208_));
 sky130_fd_sc_hs__ha_1 _11624_ (.A(\mel_ptr[0] ),
    .B(\mel_ptr[1] ),
    .COUT(_00209_),
    .SUM(_05860_));
 sky130_fd_sc_hs__ha_1 _11625_ (.A(net3609),
    .B(net3631),
    .COUT(_00212_),
    .SUM(_00213_));
 sky130_fd_sc_hs__ha_1 _11626_ (.A(net3609),
    .B(net3631),
    .COUT(_00214_),
    .SUM(_05861_));
 sky130_fd_sc_hs__ha_1 _11627_ (.A(net3608),
    .B(_00215_),
    .COUT(_00216_),
    .SUM(_00217_));
 sky130_fd_sc_hs__ha_1 _11628_ (.A(net3749),
    .B(net3748),
    .COUT(_00218_),
    .SUM(_00219_));
 sky130_fd_sc_hs__ha_1 _11629_ (.A(net3749),
    .B(net3748),
    .COUT(_00220_),
    .SUM(_05862_));
 sky130_fd_sc_hs__ha_1 _11630_ (.A(_00221_),
    .B(_00222_),
    .COUT(_00223_),
    .SUM(_00224_));
 sky130_fd_sc_hs__ha_1 _11631_ (.A(\u_window_buffer.move_counter[0] ),
    .B(_00222_),
    .COUT(_00225_),
    .SUM(_05863_));
 sky130_fd_sc_hs__ha_1 _11632_ (.A(\u_window_buffer.read_ptr[0] ),
    .B(\u_window_buffer.read_ptr[1] ),
    .COUT(_00226_),
    .SUM(_00227_));
 sky130_fd_sc_hs__ha_2 _11633_ (.A(\u_window_buffer.write_ptr[0] ),
    .B(\u_window_buffer.write_ptr[1] ),
    .COUT(_00228_),
    .SUM(_00229_));
 sky130_fd_sc_hs__ha_1 _11634_ (.A(_00230_),
    .B(_00231_),
    .COUT(_00232_),
    .SUM(_00233_));
 sky130_fd_sc_hs__ha_1 _11635_ (.A(\tx_fifo.read_ptr[0] ),
    .B(\tx_fifo.read_ptr[1] ),
    .COUT(_00234_),
    .SUM(_05864_));
 sky130_fd_sc_hs__ha_1 _11636_ (.A(_00235_),
    .B(_00236_),
    .COUT(_00237_),
    .SUM(_00238_));
 sky130_fd_sc_hs__ha_1 _11637_ (.A(\u_hamming_window.calc_pointer[0] ),
    .B(\u_hamming_window.calc_pointer[1] ),
    .COUT(_00239_),
    .SUM(_05865_));
 sky130_fd_sc_hs__ha_1 _11638_ (.A(\u_mel.k_next[0] ),
    .B(_00240_),
    .COUT(_00241_),
    .SUM(\u_mel.k_next[1] ));
 sky130_fd_sc_hs__ha_1 _11639_ (.A(\u_mel.k[0] ),
    .B(\u_mel.k[1] ),
    .COUT(_00242_),
    .SUM(_05866_));
 sky130_fd_sc_hs__dfxtp_1 _11640_ (.D(_00023_),
    .Q(_00556_),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hs__dfxtp_1 _11641_ (.D(_00024_),
    .Q(_00557_),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hs__buf_1 place2089 (.A(_04637_),
    .X(net2089));
 sky130_fd_sc_hs__buf_1 place2099 (.A(net2098),
    .X(net2099));
 sky130_fd_sc_hs__buf_1 place2087 (.A(net5133),
    .X(net2087));
 sky130_fd_sc_hs__bufbuf_8 place2088 (.A(_01791_),
    .X(net2088));
 sky130_fd_sc_hs__buf_1 place2084 (.A(net5128),
    .X(net2084));
 sky130_fd_sc_hs__buf_2 place2082 (.A(_03532_),
    .X(net2082));
 sky130_fd_sc_hs__buf_1 place2081 (.A(_03550_),
    .X(net2081));
 sky130_fd_sc_hs__buf_1 place2078 (.A(_05516_),
    .X(net2078));
 sky130_fd_sc_hs__buf_1 place2079 (.A(_04631_),
    .X(net2079));
 sky130_fd_sc_hs__buf_2 place2075 (.A(_05519_),
    .X(net2075));
 sky130_fd_sc_hs__buf_1 place2073 (.A(_03527_),
    .X(net2073));
 sky130_fd_sc_hs__buf_1 place2072 (.A(_03530_),
    .X(net2072));
 sky130_fd_sc_hs__bufbuf_8 place2071 (.A(_04633_),
    .X(net2071));
 sky130_fd_sc_hs__buf_1 place2069 (.A(net5043),
    .X(net2069));
 sky130_fd_sc_hs__buf_1 place2068 (.A(_01769_),
    .X(net2068));
 sky130_fd_sc_hs__buf_1 place2067 (.A(_01800_),
    .X(net2067));
 sky130_fd_sc_hs__bufbuf_8 place2066 (.A(_03560_),
    .X(net2066));
 sky130_fd_sc_hs__buf_1 place2065 (.A(_03563_),
    .X(net2065));
 sky130_fd_sc_hs__buf_1 place2063 (.A(_04646_),
    .X(net2063));
 sky130_fd_sc_hs__buf_1 place2062 (.A(_05523_),
    .X(net2062));
 sky130_fd_sc_hs__buf_1 place2061 (.A(_05536_),
    .X(net2061));
 sky130_fd_sc_hs__bufbuf_8 place2060 (.A(_05543_),
    .X(net2060));
 sky130_fd_sc_hs__buf_1 place2059 (.A(_05554_),
    .X(net2059));
 sky130_fd_sc_hs__buf_1 place2058 (.A(_01776_),
    .X(net2058));
 sky130_fd_sc_hs__buf_1 place2057 (.A(_01796_),
    .X(net2057));
 sky130_fd_sc_hs__buf_4 place2056 (.A(_01801_),
    .X(net2056));
 sky130_fd_sc_hs__buf_1 place2055 (.A(_01826_),
    .X(net2055));
 sky130_fd_sc_hs__buf_1 place2054 (.A(_04642_),
    .X(net2054));
 sky130_fd_sc_hs__buf_1 place2053 (.A(_04663_),
    .X(net2053));
 sky130_fd_sc_hs__buf_1 place2049 (.A(_05545_),
    .X(net2049));
 sky130_fd_sc_hs__buf_1 place2048 (.A(_01804_),
    .X(net2048));
 sky130_fd_sc_hs__buf_1 place2047 (.A(_03573_),
    .X(net2047));
 sky130_fd_sc_hs__buf_1 place2046 (.A(_03579_),
    .X(net2046));
 sky130_fd_sc_hs__buf_1 place2044 (.A(_04650_),
    .X(net2044));
 sky130_fd_sc_hs__buf_1 place2043 (.A(_05548_),
    .X(net2043));
 sky130_fd_sc_hs__buf_1 place2042 (.A(_05550_),
    .X(net2042));
 sky130_fd_sc_hs__buf_1 place2041 (.A(_01802_),
    .X(net2041));
 sky130_fd_sc_hs__buf_1 place2040 (.A(net3837),
    .X(net2040));
 sky130_fd_sc_hs__buf_1 place2045 (.A(_04644_),
    .X(net2045));
 sky130_fd_sc_hs__buf_1 place2038 (.A(_01821_),
    .X(net2038));
 sky130_fd_sc_hs__buf_1 place2037 (.A(_01864_),
    .X(net2037));
 sky130_fd_sc_hs__buf_1 place2036 (.A(_03572_),
    .X(net2036));
 sky130_fd_sc_hs__buf_1 place2035 (.A(_04647_),
    .X(net2035));
 sky130_fd_sc_hs__buf_1 place2034 (.A(_04676_),
    .X(net2034));
 sky130_fd_sc_hs__buf_1 place2029 (.A(_05579_),
    .X(net2029));
 sky130_fd_sc_hs__buf_1 place2028 (.A(_01805_),
    .X(net2028));
 sky130_fd_sc_hs__buf_2 place2026 (.A(_01836_),
    .X(net2026));
 sky130_fd_sc_hs__buf_1 place2025 (.A(_01846_),
    .X(net2025));
 sky130_fd_sc_hs__buf_1 place2027 (.A(net2026),
    .X(net2027));
 sky130_fd_sc_hs__buf_1 place2024 (.A(_03570_),
    .X(net2024));
 sky130_fd_sc_hs__buf_2 place2023 (.A(_03577_),
    .X(net2023));
 sky130_fd_sc_hs__buf_1 place2022 (.A(_03591_),
    .X(net2022));
 sky130_fd_sc_hs__buf_1 place2021 (.A(_04675_),
    .X(net2021));
 sky130_fd_sc_hs__buf_1 place2020 (.A(_05567_),
    .X(net2020));
 sky130_fd_sc_hs__bufbuf_8 place2019 (.A(_05575_),
    .X(net2019));
 sky130_fd_sc_hs__buf_1 place2018 (.A(net5091),
    .X(net2018));
 sky130_fd_sc_hs__buf_1 place2030 (.A(_05579_),
    .X(net2030));
 sky130_fd_sc_hs__buf_1 place2015 (.A(_01811_),
    .X(net2015));
 sky130_fd_sc_hs__buf_2 place2014 (.A(_01831_),
    .X(net2014));
 sky130_fd_sc_hs__buf_1 place2013 (.A(_01837_),
    .X(net2013));
 sky130_fd_sc_hs__buf_1 place2011 (.A(_03596_),
    .X(net2011));
 sky130_fd_sc_hs__bufbuf_8 place2010 (.A(_03597_),
    .X(net2010));
 sky130_fd_sc_hs__bufbuf_8 place2012 (.A(_01847_),
    .X(net2012));
 sky130_fd_sc_hs__bufbuf_8 place2009 (.A(_04658_),
    .X(net2009));
 sky130_fd_sc_hs__buf_1 place2008 (.A(_04673_),
    .X(net2008));
 sky130_fd_sc_hs__buf_1 place2007 (.A(_04679_),
    .X(net2007));
 sky130_fd_sc_hs__buf_1 place2006 (.A(_04694_),
    .X(net2006));
 sky130_fd_sc_hs__buf_1 place2005 (.A(_05588_),
    .X(net2005));
 sky130_fd_sc_hs__buf_1 place2004 (.A(net5109),
    .X(net2004));
 sky130_fd_sc_hs__buf_1 place2002 (.A(_04674_),
    .X(net2002));
 sky130_fd_sc_hs__buf_1 place2001 (.A(_04682_),
    .X(net2001));
 sky130_fd_sc_hs__buf_1 place2000 (.A(_05577_),
    .X(net2000));
 sky130_fd_sc_hs__buf_2 place1999 (.A(_03588_),
    .X(net1999));
 sky130_fd_sc_hs__buf_1 place2003 (.A(_04656_),
    .X(net2003));
 sky130_fd_sc_hs__buf_2 place1998 (.A(_04685_),
    .X(net1998));
 sky130_fd_sc_hs__buf_1 place1994 (.A(_04688_),
    .X(net1994));
 sky130_fd_sc_hs__buf_1 place1993 (.A(net5100),
    .X(net1993));
 sky130_fd_sc_hs__buf_1 place1992 (.A(_05582_),
    .X(net1992));
 sky130_fd_sc_hs__buf_1 place1995 (.A(_04688_),
    .X(net1995));
 sky130_fd_sc_hs__buf_1 place1990 (.A(_01841_),
    .X(net1990));
 sky130_fd_sc_hs__buf_1 place1991 (.A(_01838_),
    .X(net1991));
 sky130_fd_sc_hs__buf_4 place1988 (.A(_03586_),
    .X(net1988));
 sky130_fd_sc_hs__buf_1 place1984 (.A(_05581_),
    .X(net1984));
 sky130_fd_sc_hs__bufbuf_8 place1983 (.A(_01870_),
    .X(net1983));
 sky130_fd_sc_hs__buf_1 place1982 (.A(_01873_),
    .X(net1982));
 sky130_fd_sc_hs__buf_1 place1981 (.A(_03593_),
    .X(net1981));
 sky130_fd_sc_hs__buf_1 place1980 (.A(_03620_),
    .X(net1980));
 sky130_fd_sc_hs__buf_1 place1978 (.A(_04684_),
    .X(net1978));
 sky130_fd_sc_hs__buf_1 place1977 (.A(_05586_),
    .X(net1977));
 sky130_fd_sc_hs__bufbuf_8 place1976 (.A(_05592_),
    .X(net1976));
 sky130_fd_sc_hs__buf_1 place1975 (.A(_05603_),
    .X(net1975));
 sky130_fd_sc_hs__buf_1 place1973 (.A(_05624_),
    .X(net1973));
 sky130_fd_sc_hs__buf_1 place1969 (.A(_01866_),
    .X(net1969));
 sky130_fd_sc_hs__buf_1 place1967 (.A(_01899_),
    .X(net1967));
 sky130_fd_sc_hs__buf_1 place1965 (.A(_04707_),
    .X(net1965));
 sky130_fd_sc_hs__bufbuf_8 place1964 (.A(_04716_),
    .X(net1964));
 sky130_fd_sc_hs__buf_1 place1962 (.A(_05604_),
    .X(net1962));
 sky130_fd_sc_hs__buf_1 place1963 (.A(_04722_),
    .X(net1963));
 sky130_fd_sc_hs__buf_1 place1960 (.A(net5062),
    .X(net1960));
 sky130_fd_sc_hs__buf_1 place1958 (.A(_03616_),
    .X(net1958));
 sky130_fd_sc_hs__buf_1 place1957 (.A(_03631_),
    .X(net1957));
 sky130_fd_sc_hs__buf_1 place1956 (.A(_04710_),
    .X(net1956));
 sky130_fd_sc_hs__buf_1 place1954 (.A(_04738_),
    .X(net1954));
 sky130_fd_sc_hs__buf_1 place1952 (.A(_05611_),
    .X(net1952));
 sky130_fd_sc_hs__buf_1 place1953 (.A(_04739_),
    .X(net1953));
 sky130_fd_sc_hs__buf_1 place1951 (.A(_05614_),
    .X(net1951));
 sky130_fd_sc_hs__buf_1 place1950 (.A(net4867),
    .X(net1950));
 sky130_fd_sc_hs__buf_1 place1948 (.A(_03610_),
    .X(net1948));
 sky130_fd_sc_hs__buf_1 place1949 (.A(_01895_),
    .X(net1949));
 sky130_fd_sc_hs__buf_1 place1947 (.A(_04740_),
    .X(net1947));
 sky130_fd_sc_hs__buf_2 place1945 (.A(_05612_),
    .X(net1945));
 sky130_fd_sc_hs__bufbuf_8 place1944 (.A(_05636_),
    .X(net1944));
 sky130_fd_sc_hs__buf_1 place1943 (.A(_05640_),
    .X(net1943));
 sky130_fd_sc_hs__buf_1 place1941 (.A(_01875_),
    .X(net1941));
 sky130_fd_sc_hs__buf_1 place1940 (.A(_01894_),
    .X(net1940));
 sky130_fd_sc_hs__buf_1 place1939 (.A(_03627_),
    .X(net1939));
 sky130_fd_sc_hs__buf_4 place1938 (.A(_03635_),
    .X(net1938));
 sky130_fd_sc_hs__buf_1 place1936 (.A(_04744_),
    .X(net1936));
 sky130_fd_sc_hs__buf_1 place1934 (.A(_05620_),
    .X(net1934));
 sky130_fd_sc_hs__buf_1 place1935 (.A(_04760_),
    .X(net1935));
 sky130_fd_sc_hs__buf_1 place1933 (.A(net5098),
    .X(net1933));
 sky130_fd_sc_hs__buf_1 place1932 (.A(_05684_),
    .X(net1932));
 sky130_fd_sc_hs__buf_1 place1937 (.A(_03664_),
    .X(net1937));
 sky130_fd_sc_hs__buf_1 place1931 (.A(net4898),
    .X(net1931));
 sky130_fd_sc_hs__buf_1 place1930 (.A(net4893),
    .X(net1930));
 sky130_fd_sc_hs__buf_1 place1929 (.A(_01904_),
    .X(net1929));
 sky130_fd_sc_hs__buf_1 place1942 (.A(_01875_),
    .X(net1942));
 sky130_fd_sc_hs__buf_1 place1928 (.A(_01910_),
    .X(net1928));
 sky130_fd_sc_hs__buf_1 place1925 (.A(_03648_),
    .X(net1925));
 sky130_fd_sc_hs__buf_1 place1924 (.A(_03665_),
    .X(net1924));
 sky130_fd_sc_hs__buf_2 place1923 (.A(_04734_),
    .X(net1923));
 sky130_fd_sc_hs__buf_1 place1922 (.A(_05638_),
    .X(net1922));
 sky130_fd_sc_hs__buf_1 place1919 (.A(_03658_),
    .X(net1919));
 sky130_fd_sc_hs__buf_1 place1917 (.A(_04755_),
    .X(net1917));
 sky130_fd_sc_hs__buf_2 place1916 (.A(_05641_),
    .X(net1916));
 sky130_fd_sc_hs__bufbuf_8 place1915 (.A(_05672_),
    .X(net1915));
 sky130_fd_sc_hs__buf_1 place1914 (.A(_01918_),
    .X(net1914));
 sky130_fd_sc_hs__buf_1 place1913 (.A(net5191),
    .X(net1913));
 sky130_fd_sc_hs__buf_2 place1911 (.A(_03657_),
    .X(net1911));
 sky130_fd_sc_hs__buf_1 place1908 (.A(_04750_),
    .X(net1908));
 sky130_fd_sc_hs__buf_1 place1907 (.A(_05659_),
    .X(net1907));
 sky130_fd_sc_hs__buf_1 place1905 (.A(_05676_),
    .X(net1905));
 sky130_fd_sc_hs__buf_1 place1903 (.A(_01906_),
    .X(net1903));
 sky130_fd_sc_hs__buf_1 place1902 (.A(_01917_),
    .X(net1902));
 sky130_fd_sc_hs__buf_2 place1901 (.A(_03655_),
    .X(net1901));
 sky130_fd_sc_hs__buf_1 place1904 (.A(net1903),
    .X(net1904));
 sky130_fd_sc_hs__buf_1 place1900 (.A(_03683_),
    .X(net1900));
 sky130_fd_sc_hs__buf_1 place1898 (.A(_04749_),
    .X(net1898));
 sky130_fd_sc_hs__buf_1 place1906 (.A(_05676_),
    .X(net1906));
 sky130_fd_sc_hs__buf_2 place1896 (.A(_04773_),
    .X(net1896));
 sky130_fd_sc_hs__buf_4 place1895 (.A(_05654_),
    .X(net1895));
 sky130_fd_sc_hs__buf_1 place1894 (.A(_05664_),
    .X(net1894));
 sky130_fd_sc_hs__buf_1 place1893 (.A(_05683_),
    .X(net1893));
 sky130_fd_sc_hs__buf_2 place1891 (.A(_01919_),
    .X(net1891));
 sky130_fd_sc_hs__buf_1 place1892 (.A(net1891),
    .X(net1892));
 sky130_fd_sc_hs__buf_1 place1897 (.A(net1896),
    .X(net1897));
 sky130_fd_sc_hs__buf_1 place1890 (.A(net4873),
    .X(net1890));
 sky130_fd_sc_hs__buf_1 place1889 (.A(_01945_),
    .X(net1889));
 sky130_fd_sc_hs__bufbuf_8 place1888 (.A(_04751_),
    .X(net1888));
 sky130_fd_sc_hs__bufbuf_8 place1887 (.A(_04759_),
    .X(net1887));
 sky130_fd_sc_hs__bufbuf_8 place1886 (.A(_04769_),
    .X(net1886));
 sky130_fd_sc_hs__bufbuf_8 place1885 (.A(_04781_),
    .X(net1885));
 sky130_fd_sc_hs__buf_1 place1884 (.A(_01935_),
    .X(net1884));
 sky130_fd_sc_hs__buf_1 place1883 (.A(net4928),
    .X(net1883));
 sky130_fd_sc_hs__buf_1 place1909 (.A(_03677_),
    .X(net1909));
 sky130_fd_sc_hs__buf_1 place1882 (.A(net4894),
    .X(net1882));
 sky130_fd_sc_hs__buf_1 place1880 (.A(_01974_),
    .X(net1880));
 sky130_fd_sc_hs__buf_1 place1881 (.A(_01974_),
    .X(net1881));
 sky130_fd_sc_hs__bufbuf_8 place1879 (.A(net4889),
    .X(net1879));
 sky130_fd_sc_hs__buf_1 place1877 (.A(_05674_),
    .X(net1877));
 sky130_fd_sc_hs__buf_1 rebuffer5107 (.A(_05677_),
    .X(net5107));
 sky130_fd_sc_hs__buf_4 place1876 (.A(_01947_),
    .X(net1876));
 sky130_fd_sc_hs__buf_16 place1875 (.A(net3787),
    .X(net1875));
 sky130_fd_sc_hs__buf_16 place1874 (.A(_03673_),
    .X(net1874));
 sky130_fd_sc_hs__buf_1 place1870 (.A(_05699_),
    .X(net1870));
 sky130_fd_sc_hs__buf_2 place1871 (.A(_04771_),
    .X(net1871));
 sky130_fd_sc_hs__buf_8 place1868 (.A(_01949_),
    .X(net1868));
 sky130_fd_sc_hs__buf_1 rebuffer5190 (.A(_03445_),
    .X(net5190));
 sky130_fd_sc_hs__buf_1 place1864 (.A(_05696_),
    .X(net1864));
 sky130_fd_sc_hs__buf_8 place1861 (.A(_00456_),
    .X(net1861));
 sky130_fd_sc_hs__buf_1 place1860 (.A(_05680_),
    .X(net1860));
 sky130_fd_sc_hs__buf_1 place1859 (.A(_05693_),
    .X(net1859));
 sky130_fd_sc_hs__buf_1 place1858 (.A(net5084),
    .X(net1858));
 sky130_fd_sc_hs__buf_8 place1857 (.A(_05700_),
    .X(net1857));
 sky130_fd_sc_hs__buf_1 place1856 (.A(_05707_),
    .X(net1856));
 sky130_fd_sc_hs__bufbuf_8 place1855 (.A(_05714_),
    .X(net1855));
 sky130_fd_sc_hs__buf_2 place1854 (.A(net5199),
    .X(net1854));
 sky130_fd_sc_hs__buf_4 place1850 (.A(_05757_),
    .X(net1850));
 sky130_fd_sc_hs__buf_8 rebuffer5262 (.A(_03686_),
    .X(net5262));
 sky130_fd_sc_hs__buf_8 place1849 (.A(_05722_),
    .X(net1849));
 sky130_fd_sc_hs__buf_8 place1848 (.A(_02119_),
    .X(net1848));
 sky130_fd_sc_hs__buf_1 place1852 (.A(_05720_),
    .X(net1852));
 sky130_fd_sc_hs__clkbuf_16 place1845 (.A(_03868_),
    .X(net1845));
 sky130_fd_sc_hs__buf_8 place1844 (.A(_02121_),
    .X(net1844));
 sky130_fd_sc_hs__buf_16 rebuffer4958 (.A(_04787_),
    .X(net4958));
 sky130_fd_sc_hs__buf_8 place1841 (.A(_02770_),
    .X(net1841));
 sky130_fd_sc_hs__buf_16 place1840 (.A(_00022_),
    .X(net1840));
 sky130_fd_sc_hs__clkbuf_16 place1846 (.A(net1845),
    .X(net1846));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hs__clkbuf_16 place1842 (.A(_04792_),
    .X(net1842));
 sky130_fd_sc_hs__buf_4 place3780 (.A(_05774_),
    .X(net3780));
 sky130_fd_sc_hs__buf_1 place3679 (.A(\u_window_buffer.write_ptr[8] ),
    .X(net3679));
 sky130_fd_sc_hs__buf_1 output213 (.A(net213),
    .X(mfcc_done_o));
 sky130_fd_sc_hs__buf_1 input212 (.A(start_i),
    .X(net212));
 sky130_fd_sc_hs__clkbuf_4 input211 (.A(rst_n),
    .X(net211));
 sky130_fd_sc_hs__buf_1 input210 (.A(pcm_ready_i),
    .X(net210));
 sky130_fd_sc_hs__buf_1 input209 (.A(auto_restart_i),
    .X(net209));
 sky130_fd_sc_hs__dfxtp_1 \hamming_finished$_SDFFE_PP0P_  (.D(_00243_),
    .Q(hamming_finished),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hs__edfxtp_1 \start_move$_DFFE_PN_  (.D(_00000_),
    .DE(_05774_),
    .Q(start_move),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hs__dfxtp_1 \start_move_auto$_SDFF_PN0_  (.D(_00244_),
    .Q(start_move_auto),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.read_ptr[0]$_SDFFE_PN0P_  (.D(_00245_),
    .Q(\tx_fifo.read_ptr[0] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.read_ptr[1]$_SDFFE_PN0P_  (.D(_00246_),
    .Q(\tx_fifo.read_ptr[1] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.read_ptr[2]$_SDFFE_PN0P_  (.D(_00247_),
    .Q(\tx_fifo.read_ptr[2] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.read_ptr[3]$_SDFFE_PN0P_  (.D(_00248_),
    .Q(\tx_fifo.read_ptr[3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.read_ptr[4]$_SDFFE_PN0P_  (.D(_00249_),
    .Q(\tx_fifo.read_ptr[4] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.read_ptr[5]$_SDFFE_PN0P_  (.D(_00250_),
    .Q(\tx_fifo.read_ptr[5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.read_ptr[6]$_SDFFE_PN0P_  (.D(_00251_),
    .Q(\tx_fifo.read_ptr[6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.read_ptr[7]$_SDFFE_PN0P_  (.D(_00252_),
    .Q(\tx_fifo.read_ptr[7] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.write_ptr[0]$_SDFFE_PN0P_  (.D(_00253_),
    .Q(\tx_fifo.write_ptr[0] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.write_ptr[1]$_SDFFE_PN0P_  (.D(_00254_),
    .Q(\tx_fifo.write_ptr[1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.write_ptr[2]$_SDFFE_PN0P_  (.D(_00255_),
    .Q(\tx_fifo.write_ptr[2] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.write_ptr[3]$_SDFFE_PN0P_  (.D(_00256_),
    .Q(\tx_fifo.write_ptr[3] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.write_ptr[4]$_SDFFE_PN0P_  (.D(_00257_),
    .Q(\tx_fifo.write_ptr[4] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.write_ptr[5]$_SDFFE_PN0P_  (.D(_00258_),
    .Q(\tx_fifo.write_ptr[5] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.write_ptr[6]$_SDFFE_PN0P_  (.D(_00259_),
    .Q(\tx_fifo.write_ptr[6] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hs__dfxtp_1 \tx_fifo.write_ptr[7]$_SDFFE_PN0P_  (.D(_00260_),
    .Q(\tx_fifo.write_ptr[7] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.dct_done_o$_SDFF_PN0_  (.D(_00261_),
    .Q(net213),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.dct_state[0]$_DFF_P_  (.D(_00007_),
    .Q(\u_dct.dct_state[0] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.dct_state[1]$_DFF_P_  (.D(_00001_),
    .Q(\u_dct.dct_state[1] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.dct_state[2]$_DFF_P_  (.D(_00008_),
    .Q(\u_dct.dct_state[2] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.dct_state[3]$_DFF_P_  (.D(_00002_),
    .Q(\u_dct.dct_state[3] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.k_ptr[0]$_SDFFE_PN0P_  (.D(_00262_),
    .Q(\u_dct.k_ptr[0] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.k_ptr[1]$_SDFFE_PN0P_  (.D(_00263_),
    .Q(\u_dct.k_ptr[1] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.k_ptr[2]$_SDFFE_PN0P_  (.D(_00264_),
    .Q(\u_dct.k_ptr[2] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.k_ptr[3]$_SDFFE_PN0P_  (.D(_00265_),
    .Q(\u_dct.k_ptr[3] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.n_ptr[0]$_SDFFE_PN0P_  (.D(_00266_),
    .Q(\u_dct.n_ptr[0] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.n_ptr[1]$_SDFFE_PN0P_  (.D(_00267_),
    .Q(\u_dct.n_ptr[1] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.n_ptr[2]$_SDFFE_PN0P_  (.D(_00268_),
    .Q(\u_dct.n_ptr[2] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.n_ptr[3]$_SDFFE_PN0P_  (.D(_00269_),
    .Q(\u_dct.n_ptr[3] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.n_ptr[4]$_SDFFE_PN0P_  (.D(_00270_),
    .Q(\u_dct.n_ptr[4] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_dct.n_ptr[5]$_SDFFE_PN0P_  (.D(_00271_),
    .Q(\u_dct.n_ptr[5] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.fft_done_o$_SDFF_PN0_  (.D(_00272_),
    .Q(fft_done),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.fft_state[0]$_DFF_P_  (.D(_00009_),
    .Q(\u_fft.fft_state[0] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.fft_state[1]$_DFF_P_  (.D(_00010_),
    .Q(\u_fft.fft_state[1] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.fft_state[2]$_DFF_P_  (.D(_00011_),
    .Q(\u_fft.fft_state[2] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.fft_state[3]$_DFF_P_  (.D(_00003_),
    .Q(\u_fft.fft_state[3] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr[0]$_SDFFE_PN0P_  (.D(_00273_),
    .Q(\u_fft.power_ptr[0] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr[1]$_SDFFE_PN0P_  (.D(_00274_),
    .Q(\u_fft.power_ptr[1] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr[2]$_SDFFE_PN0P_  (.D(_00275_),
    .Q(\u_fft.power_ptr[2] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr[3]$_SDFFE_PN0P_  (.D(_00276_),
    .Q(\u_fft.power_ptr[3] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr[4]$_SDFFE_PN0P_  (.D(_00277_),
    .Q(\u_fft.power_ptr[4] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr[5]$_SDFFE_PN0P_  (.D(_00278_),
    .Q(\u_fft.power_ptr[5] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr[6]$_SDFFE_PN0P_  (.D(_00279_),
    .Q(\u_fft.power_ptr[6] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr[7]$_SDFFE_PN0P_  (.D(_00280_),
    .Q(\u_fft.power_ptr[7] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr[8]$_SDFFE_PN0P_  (.D(_00281_),
    .Q(\u_fft.power_ptr[8] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr[9]$_SDFFE_PN0P_  (.D(_00282_),
    .Q(\u_fft.power_ptr[9] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage1[0]$_SDFFE_PN0P_  (.D(_00283_),
    .Q(\u_fft.power_ptr_stage1[0] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage1[1]$_SDFFE_PN0P_  (.D(_00284_),
    .Q(\u_fft.power_ptr_stage1[1] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage1[2]$_SDFFE_PN0P_  (.D(_00285_),
    .Q(\u_fft.power_ptr_stage1[2] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage1[3]$_SDFFE_PN0P_  (.D(_00286_),
    .Q(\u_fft.power_ptr_stage1[3] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage1[4]$_SDFFE_PN0P_  (.D(_00287_),
    .Q(\u_fft.power_ptr_stage1[4] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage1[5]$_SDFFE_PN0P_  (.D(_00288_),
    .Q(\u_fft.power_ptr_stage1[5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage1[6]$_SDFFE_PN0P_  (.D(_00289_),
    .Q(\u_fft.power_ptr_stage1[6] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage1[7]$_SDFFE_PN0P_  (.D(_00290_),
    .Q(\u_fft.power_ptr_stage1[7] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage1[8]$_SDFFE_PN0P_  (.D(_00291_),
    .Q(\u_fft.power_ptr_stage1[8] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage1[9]$_SDFFE_PN0P_  (.D(_00292_),
    .Q(\u_fft.power_ptr_stage1[9] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage2[0]$_SDFFE_PN0P_  (.D(_00293_),
    .Q(\u_fft.power_ptr_stage2[0] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage2[1]$_SDFFE_PN0P_  (.D(_00294_),
    .Q(\u_fft.power_ptr_stage2[1] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage2[2]$_SDFFE_PN0P_  (.D(_00295_),
    .Q(\u_fft.power_ptr_stage2[2] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage2[3]$_SDFFE_PN0P_  (.D(_00296_),
    .Q(\u_fft.power_ptr_stage2[3] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage2[4]$_SDFFE_PN0P_  (.D(_00297_),
    .Q(\u_fft.power_ptr_stage2[4] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage2[5]$_SDFFE_PN0P_  (.D(_00298_),
    .Q(\u_fft.power_ptr_stage2[5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage2[6]$_SDFFE_PN0P_  (.D(_00299_),
    .Q(\u_fft.power_ptr_stage2[6] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage2[7]$_SDFFE_PN0P_  (.D(_00300_),
    .Q(\u_fft.power_ptr_stage2[7] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage2[8]$_SDFFE_PN0P_  (.D(_00301_),
    .Q(\u_fft.power_ptr_stage2[8] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage2[9]$_SDFFE_PN0P_  (.D(_00302_),
    .Q(\u_fft.power_ptr_stage2[9] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage3[0]$_SDFFE_PN0P_  (.D(_00303_),
    .Q(\u_fft.power_ptr_stage3[0] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage3[1]$_SDFFE_PN0P_  (.D(_00304_),
    .Q(\u_fft.power_ptr_stage3[1] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage3[2]$_SDFFE_PN0P_  (.D(_00305_),
    .Q(\u_fft.power_ptr_stage3[2] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage3[3]$_SDFFE_PN0P_  (.D(_00306_),
    .Q(\u_fft.power_ptr_stage3[3] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage3[4]$_SDFFE_PN0P_  (.D(_00307_),
    .Q(\u_fft.power_ptr_stage3[4] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage3[5]$_SDFFE_PN0P_  (.D(_00308_),
    .Q(\u_fft.power_ptr_stage3[5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage3[6]$_SDFFE_PN0P_  (.D(_00309_),
    .Q(\u_fft.power_ptr_stage3[6] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage3[7]$_SDFFE_PN0P_  (.D(_00310_),
    .Q(\u_fft.power_ptr_stage3[7] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage3[8]$_SDFFE_PN0P_  (.D(_00311_),
    .Q(\u_fft.power_ptr_stage3[8] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage3[9]$_SDFFE_PN0P_  (.D(_00312_),
    .Q(\u_fft.power_ptr_stage3[9] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage4[0]$_SDFFE_PN0P_  (.D(_00313_),
    .Q(\fft_ptr[0] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage4[1]$_SDFFE_PN0P_  (.D(_00314_),
    .Q(\fft_ptr[1] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage4[2]$_SDFFE_PN0P_  (.D(_00315_),
    .Q(\fft_ptr[2] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage4[3]$_SDFFE_PN0P_  (.D(_00316_),
    .Q(\fft_ptr[3] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage4[4]$_SDFFE_PN0P_  (.D(_00317_),
    .Q(\fft_ptr[4] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage4[5]$_SDFFE_PN0P_  (.D(_00318_),
    .Q(\fft_ptr[5] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage4[6]$_SDFFE_PN0P_  (.D(_00319_),
    .Q(\fft_ptr[6] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage4[7]$_SDFFE_PN0P_  (.D(_00320_),
    .Q(\fft_ptr[7] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage4[8]$_SDFFE_PN0P_  (.D(_00321_),
    .Q(\fft_ptr[8] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.power_ptr_stage4[9]$_SDFFE_PN0P_  (.D(_00322_),
    .Q(\u_fft.power_ptr_stage4[9] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[20]$_SDFFE_PN1P_  (.D(_00323_),
    .Q(\u_fft.sched[20] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[21]$_SDFFE_PN0P_  (.D(_00324_),
    .Q(\u_fft.sched[21] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[22]$_SDFFE_PN0P_  (.D(_00325_),
    .Q(\u_fft.sched[22] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[23]$_SDFFE_PN0P_  (.D(_00326_),
    .Q(\u_fft.sched[23] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[24]$_SDFFE_PN0P_  (.D(_00327_),
    .Q(\u_fft.sched[24] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[25]$_SDFFE_PN0P_  (.D(_00328_),
    .Q(\u_fft.sched[25] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[26]$_SDFFE_PN0P_  (.D(_00329_),
    .Q(\u_fft.sched[26] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[27]$_SDFFE_PN0P_  (.D(_00330_),
    .Q(\u_fft.sched[1] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[28]$_SDFFE_PN0P_  (.D(_00331_),
    .Q(\u_fft.sched[0] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[29]$_SDFFE_PN0P_  (.D(_00332_),
    .Q(\u_fft.sched[29] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[30]$_SDFFE_PN0P_  (.D(_00333_),
    .Q(\u_fft.sched[30] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[31]$_SDFFE_PN1P_  (.D(_00334_),
    .Q(\u_fft.sched[31] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[32]$_SDFFE_PN0P_  (.D(_00335_),
    .Q(\u_fft.sched[32] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[33]$_SDFFE_PN0P_  (.D(_00336_),
    .Q(\u_fft.sched[33] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[34]$_SDFFE_PN0P_  (.D(_00337_),
    .Q(\u_fft.sched[34] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[35]$_SDFFE_PN0P_  (.D(_00338_),
    .Q(\u_fft.sched[35] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[36]$_SDFFE_PN0P_  (.D(_00339_),
    .Q(\u_fft.sched[36] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[37]$_SDFFE_PN0P_  (.D(_00340_),
    .Q(\u_fft.sched[37] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[38]$_SDFFE_PN0P_  (.D(_00341_),
    .Q(\u_fft.sched[38] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[39]$_SDFFE_PN0P_  (.D(_00342_),
    .Q(\u_fft.sched[39] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[40]$_SDFFE_PN1P_  (.D(_00343_),
    .Q(\u_fft.sched[40] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[41]$_SDFFE_PN0P_  (.D(_00344_),
    .Q(\u_fft.sched[41] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[42]$_SDFFE_PN0P_  (.D(_00345_),
    .Q(\u_fft.sched[42] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[43]$_SDFFE_PN0P_  (.D(_00346_),
    .Q(\u_fft.sched[43] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[44]$_SDFFE_PN0P_  (.D(_00347_),
    .Q(\u_fft.sched[44] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[45]$_SDFFE_PN0P_  (.D(_00348_),
    .Q(\u_fft.sched[45] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[46]$_SDFFE_PN0P_  (.D(_00349_),
    .Q(\u_fft.sched[46] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[47]$_SDFFE_PN0P_  (.D(_00350_),
    .Q(\u_fft.sched[47] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[48]$_SDFFE_PN0P_  (.D(_00351_),
    .Q(\u_fft.sched[48] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[49]$_SDFFE_PN0P_  (.D(_00352_),
    .Q(\u_fft.sched[49] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[50]$_SDFFE_PN0P_  (.D(_00353_),
    .Q(\u_fft.sched[50] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[51]$_SDFFE_PN0P_  (.D(_00354_),
    .Q(\u_fft.sched[51] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[52]$_SDFFE_PN0P_  (.D(_00355_),
    .Q(\u_fft.sched[52] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[53]$_SDFFE_PN0P_  (.D(_00356_),
    .Q(\u_fft.sched[53] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[54]$_SDFFE_PN0P_  (.D(_00357_),
    .Q(\u_fft.sched[54] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[55]$_SDFFE_PN0P_  (.D(_00358_),
    .Q(\u_fft.sched[55] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[56]$_SDFFE_PN0P_  (.D(_00359_),
    .Q(\u_fft.sched[56] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[57]$_SDFFE_PN0P_  (.D(_00360_),
    .Q(\u_fft.sched[57] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[58]$_SDFFE_PN0P_  (.D(_00361_),
    .Q(\u_fft.sched[58] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[59]$_SDFFE_PN0P_  (.D(_00362_),
    .Q(\u_fft.sched[59] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[60]$_SDFFE_PN0P_  (.D(_00363_),
    .Q(\u_fft.sched[60] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[61]$_SDFFE_PN0P_  (.D(_00364_),
    .Q(\u_fft.sched[61] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[62]$_SDFFE_PN0P_  (.D(_00365_),
    .Q(\u_fft.sched[62] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[63]$_SDFFE_PN0P_  (.D(_00366_),
    .Q(\u_fft.sched[63] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_fft.sched[64]$_SDFFE_PN0P_  (.D(_00367_),
    .Q(\u_fft.sched[64] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[0]$_SDFFCE_PN0P_  (.D(_00368_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[0] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[10]$_SDFFCE_PN0P_  (.D(_00369_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[10] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[11]$_SDFFCE_PN0P_  (.D(_00370_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[11] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[12]$_SDFFCE_PN0P_  (.D(_00371_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[12] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[13]$_SDFFCE_PN0P_  (.D(_00372_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[13] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[14]$_SDFFCE_PN0P_  (.D(_00373_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[14] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[15]$_SDFFCE_PN0P_  (.D(_00374_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[15] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[16]$_SDFFCE_PN0P_  (.D(_00375_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[16] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[17]$_SDFFCE_PN0P_  (.D(_00376_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[17] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[18]$_SDFFCE_PN0P_  (.D(_00377_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[18] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[19]$_SDFFCE_PN0P_  (.D(_00378_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[19] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[1]$_SDFFCE_PN0P_  (.D(_00379_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[1] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[20]$_SDFFCE_PN0P_  (.D(_00380_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[20] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[21]$_SDFFCE_PN0P_  (.D(_00381_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[21] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[22]$_SDFFCE_PN0P_  (.D(_00382_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[22] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[23]$_SDFFCE_PN0P_  (.D(_00383_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[23] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[24]$_SDFFCE_PN0P_  (.D(_00384_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[24] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[25]$_SDFFCE_PN0P_  (.D(_00385_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[25] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[26]$_SDFFCE_PN0P_  (.D(_00386_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[26] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[27]$_SDFFCE_PN0P_  (.D(_00387_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[27] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[28]$_SDFFCE_PN0P_  (.D(_00388_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[28] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[29]$_SDFFCE_PN0P_  (.D(_00389_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[29] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[2]$_SDFFCE_PN0P_  (.D(_00390_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[2] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[30]$_SDFFCE_PN0P_  (.D(_00391_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[31]$_SDFFCE_PN0P_  (.D(_00392_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[31] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[3]$_SDFFCE_PN0P_  (.D(_00393_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[3] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[4]$_SDFFCE_PN0P_  (.D(_00394_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[4] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[5]$_SDFFCE_PN0P_  (.D(_00395_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[5] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[6]$_SDFFCE_PN0P_  (.D(_00396_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[6] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[7]$_SDFFCE_PN0P_  (.D(_00397_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[7] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[8]$_SDFFCE_PN0P_  (.D(_00398_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[8] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_hamming_window.calc_pointer[9]$_SDFFCE_PN0P_  (.D(_00399_),
    .DE(net1840),
    .Q(\u_hamming_window.calc_pointer[9] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.done$_SDFF_PN0_  (.D(_00400_),
    .Q(\u_hamming_window.done ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.done_o$_DFF_P_  (.D(\u_hamming_window.done ),
    .Q(hamming_done),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.frame_ptr[0]$_SDFFE_PN0P_  (.D(_00401_),
    .Q(\u_hamming_window.frame_ptr[0] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.frame_ptr[1]$_SDFFE_PN0P_  (.D(_00402_),
    .Q(\u_hamming_window.frame_ptr[1] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.frame_ptr[2]$_SDFFE_PN0P_  (.D(_00403_),
    .Q(\u_hamming_window.frame_ptr[2] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.frame_ptr[3]$_SDFFE_PN0P_  (.D(_00404_),
    .Q(\u_hamming_window.frame_ptr[3] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.frame_ptr[4]$_SDFFE_PN0P_  (.D(_00405_),
    .Q(\u_hamming_window.frame_ptr[4] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.frame_ptr[5]$_SDFFE_PN0P_  (.D(_00406_),
    .Q(\u_hamming_window.frame_ptr[5] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.frame_ptr[6]$_SDFFE_PN0P_  (.D(_00407_),
    .Q(\u_hamming_window.frame_ptr[6] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.frame_ptr[7]$_SDFFE_PN0P_  (.D(_00408_),
    .Q(\u_hamming_window.frame_ptr[7] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.frame_ptr[8]$_SDFFE_PN0P_  (.D(_00409_),
    .Q(\u_hamming_window.frame_ptr[8] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.hamming_state[0]$_DFF_P_  (.D(_00012_),
    .Q(\u_hamming_window.hamming_state[0] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.hamming_state[1]$_DFF_P_  (.D(_00013_),
    .Q(\u_hamming_window.hamming_state[1] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.hamming_state[2]$_DFF_P_  (.D(_00014_),
    .Q(\u_hamming_window.hamming_state[2] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.hamming_state[3]$_DFF_P_  (.D(_00004_),
    .Q(\u_hamming_window.hamming_state[3] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_hamming_window.rd_en_o$_SDFF_PN0_  (.D(_00410_),
    .Q(\u_hamming_window.rd_en_o ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.k[0]$_SDFFE_PN0P_  (.D(_00411_),
    .Q(\u_mel.k[0] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.k[1]$_SDFFE_PN0P_  (.D(_00412_),
    .Q(\u_mel.k[1] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.k[2]$_SDFFE_PN0P_  (.D(_00413_),
    .Q(\u_mel.k[2] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.k[3]$_SDFFE_PN0P_  (.D(_00414_),
    .Q(\u_mel.k[3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.k[4]$_SDFFE_PN0P_  (.D(_00415_),
    .Q(\u_mel.k[4] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.k[5]$_SDFFE_PN0P_  (.D(_00416_),
    .Q(\u_mel.k[5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.k[6]$_SDFFE_PN0P_  (.D(_00417_),
    .Q(\u_mel.k[6] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.k[7]$_SDFFE_PN0P_  (.D(_00418_),
    .Q(\u_mel.k[7] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.k[8]$_SDFFE_PN0P_  (.D(_00419_),
    .Q(\u_mel.k[8] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.mel_done_o$_SDFF_PN0_  (.D(_00420_),
    .Q(mel_done),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.mel_prt_energies[0]$_SDFFE_PN0P_  (.D(_00421_),
    .Q(\mel_ptr[0] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.mel_prt_energies[1]$_SDFFE_PN0P_  (.D(_00422_),
    .Q(\mel_ptr[1] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.mel_prt_energies[2]$_SDFFE_PN0P_  (.D(_00423_),
    .Q(\mel_ptr[2] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.mel_prt_energies[3]$_SDFFE_PN0P_  (.D(_00424_),
    .Q(\mel_ptr[3] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.mel_prt_energies[4]$_SDFFE_PN0P_  (.D(_00425_),
    .Q(\mel_ptr[4] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.mel_prt_energies[5]$_SDFFE_PN0P_  (.D(_00426_),
    .Q(\mel_ptr[5] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.state[0]$_DFF_P_  (.D(_00015_),
    .Q(\u_mel.state[0] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.state[1]$_DFF_P_  (.D(_00016_),
    .Q(\u_mel.state[1] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.state[2]$_DFF_P_  (.D(_00017_),
    .Q(\u_mel.state[2] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_mel.state[3]$_DFF_P_  (.D(_00005_),
    .Q(mel_valid),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hs__edfxtp_1 \u_pre_emphasis.out_valid$_DFFE_PP_  (.D(net210),
    .DE(net211),
    .Q(pre_emphasis_valid),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.current_state[0]$_DFF_P_  (.D(net3782),
    .Q(\u_window_buffer.current_state[0] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.current_state[1]$_DFF_P_  (.D(_00019_),
    .Q(idle),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.current_state[2]$_DFF_P_  (.D(_00020_),
    .Q(\u_window_buffer.current_state[2] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.current_state[3]$_DFF_P_  (.D(_00006_),
    .Q(\u_window_buffer.current_state[3] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.current_state[4]$_DFF_P_  (.D(_00021_),
    .Q(\u_window_buffer.current_state[4] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.fifo_rd_en_o$_SDFF_PN0_  (.D(_00427_),
    .Q(fifo_rd_en),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hs__dfxtp_4 \u_window_buffer.internal_read_ptr[10]$_SDFFE_PN0N_  (.D(_00428_),
    .Q(\u_window_buffer.internal_read_ptr[10] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hs__dfxtp_4 \u_window_buffer.internal_read_ptr[11]$_SDFFE_PN0N_  (.D(_00429_),
    .Q(\u_window_buffer.internal_read_ptr[11] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.internal_read_ptr[12]$_SDFFE_PN0N_  (.D(_00430_),
    .Q(\u_window_buffer.internal_read_ptr[12] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[13]$_SDFFE_PN0N_  (.D(_00431_),
    .Q(\u_window_buffer.internal_read_ptr[13] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hs__dfxtp_4 \u_window_buffer.internal_read_ptr[14]$_SDFFE_PN0N_  (.D(_00432_),
    .Q(\u_window_buffer.internal_read_ptr[14] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.internal_read_ptr[15]$_SDFFE_PN0N_  (.D(_00433_),
    .Q(\u_window_buffer.internal_read_ptr[15] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[16]$_SDFFE_PN0N_  (.D(_00434_),
    .Q(\u_window_buffer.internal_read_ptr[16] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.internal_read_ptr[17]$_SDFFE_PN0N_  (.D(_00435_),
    .Q(\u_window_buffer.internal_read_ptr[17] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[18]$_SDFFE_PN0N_  (.D(_00436_),
    .Q(\u_window_buffer.internal_read_ptr[18] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[19]$_SDFFE_PN0N_  (.D(_00437_),
    .Q(\u_window_buffer.internal_read_ptr[19] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[1]$_SDFFE_PN0N_  (.D(_00438_),
    .Q(\u_window_buffer.internal_read_ptr[1] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.internal_read_ptr[20]$_SDFFE_PN0N_  (.D(_00439_),
    .Q(\u_window_buffer.internal_read_ptr[20] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.internal_read_ptr[21]$_SDFFE_PN0N_  (.D(_00440_),
    .Q(\u_window_buffer.internal_read_ptr[21] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[22]$_SDFFE_PN0N_  (.D(_00441_),
    .Q(\u_window_buffer.internal_read_ptr[22] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[23]$_SDFFE_PN0N_  (.D(_00442_),
    .Q(\u_window_buffer.internal_read_ptr[23] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[24]$_SDFFE_PN0N_  (.D(_00443_),
    .Q(\u_window_buffer.internal_read_ptr[24] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[25]$_SDFFE_PN0N_  (.D(_00444_),
    .Q(\u_window_buffer.internal_read_ptr[25] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[26]$_SDFFE_PN0N_  (.D(_00445_),
    .Q(\u_window_buffer.internal_read_ptr[26] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[27]$_SDFFE_PN0N_  (.D(_00446_),
    .Q(\u_window_buffer.internal_read_ptr[27] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[28]$_SDFFE_PN0N_  (.D(_00447_),
    .Q(\u_window_buffer.internal_read_ptr[28] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[29]$_SDFFE_PN0N_  (.D(_00448_),
    .Q(\u_window_buffer.internal_read_ptr[29] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hs__dfxtp_4 \u_window_buffer.internal_read_ptr[2]$_SDFFE_PN0N_  (.D(_00449_),
    .Q(\u_window_buffer.internal_read_ptr[2] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[30]$_SDFFE_PN0N_  (.D(_00450_),
    .Q(\u_window_buffer.internal_read_ptr[30] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[31]$_SDFFE_PN0N_  (.D(_00451_),
    .Q(\u_window_buffer.internal_read_ptr[31] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hs__dfxtp_4 \u_window_buffer.internal_read_ptr[3]$_SDFFE_PN0N_  (.D(_00452_),
    .Q(\u_window_buffer.internal_read_ptr[3] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[4]$_SDFFE_PN0N_  (.D(_00453_),
    .Q(\u_window_buffer.internal_read_ptr[4] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hs__dfxtp_4 \u_window_buffer.internal_read_ptr[5]$_SDFFE_PN0N_  (.D(_00454_),
    .Q(\u_window_buffer.internal_read_ptr[5] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.internal_read_ptr[6]$_SDFFE_PN0N_  (.D(_00455_),
    .Q(\u_window_buffer.internal_read_ptr[6] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[7]$_SDFFE_PN0N_  (.D(net1861),
    .Q(\u_window_buffer.internal_read_ptr[7] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.internal_read_ptr[8]$_SDFFE_PN0N_  (.D(_00457_),
    .Q(\u_window_buffer.internal_read_ptr[8] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hs__dfxtp_4 \u_window_buffer.internal_read_ptr[9]$_SDFFE_PN0N_  (.D(_00458_),
    .Q(\u_window_buffer.internal_read_ptr[9] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[0]$_SDFFE_PN0P_  (.D(_00459_),
    .Q(\u_window_buffer.move_counter[0] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[10]$_SDFFE_PN0P_  (.D(_00460_),
    .Q(\u_window_buffer.move_counter[10] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[11]$_SDFFE_PN0P_  (.D(_00461_),
    .Q(\u_window_buffer.move_counter[11] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[12]$_SDFFE_PN0P_  (.D(_00462_),
    .Q(\u_window_buffer.move_counter[12] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[13]$_SDFFE_PN0P_  (.D(_00463_),
    .Q(\u_window_buffer.move_counter[13] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[14]$_SDFFE_PN0P_  (.D(_00464_),
    .Q(\u_window_buffer.move_counter[14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[15]$_SDFFE_PN0P_  (.D(_00465_),
    .Q(\u_window_buffer.move_counter[15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[16]$_SDFFE_PN0P_  (.D(_00466_),
    .Q(\u_window_buffer.move_counter[16] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[17]$_SDFFE_PN0P_  (.D(_00467_),
    .Q(\u_window_buffer.move_counter[17] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[18]$_SDFFE_PN0P_  (.D(_00468_),
    .Q(\u_window_buffer.move_counter[18] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[19]$_SDFFE_PN0P_  (.D(_00469_),
    .Q(\u_window_buffer.move_counter[19] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[1]$_SDFFE_PN0P_  (.D(_00470_),
    .Q(\u_window_buffer.move_counter[1] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[20]$_SDFFE_PN0P_  (.D(_00471_),
    .Q(\u_window_buffer.move_counter[20] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[21]$_SDFFE_PN0P_  (.D(_00472_),
    .Q(\u_window_buffer.move_counter[21] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[22]$_SDFFE_PN0P_  (.D(_00473_),
    .Q(\u_window_buffer.move_counter[22] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[23]$_SDFFE_PN0P_  (.D(_00474_),
    .Q(\u_window_buffer.move_counter[23] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[24]$_SDFFE_PN0P_  (.D(_00475_),
    .Q(\u_window_buffer.move_counter[24] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[25]$_SDFFE_PN0P_  (.D(_00476_),
    .Q(\u_window_buffer.move_counter[25] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[26]$_SDFFE_PN0P_  (.D(_00477_),
    .Q(\u_window_buffer.move_counter[26] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[27]$_SDFFE_PN0P_  (.D(_00478_),
    .Q(\u_window_buffer.move_counter[27] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[28]$_SDFFE_PN0P_  (.D(_00479_),
    .Q(\u_window_buffer.move_counter[28] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[29]$_SDFFE_PN0P_  (.D(_00480_),
    .Q(\u_window_buffer.move_counter[29] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[2]$_SDFFE_PN0P_  (.D(_00481_),
    .Q(\u_window_buffer.move_counter[2] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[30]$_SDFFE_PN0P_  (.D(_00482_),
    .Q(\u_window_buffer.move_counter[30] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[31]$_SDFFE_PN0P_  (.D(_00483_),
    .Q(\u_window_buffer.move_counter[31] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[3]$_SDFFE_PN0P_  (.D(_00484_),
    .Q(\u_window_buffer.move_counter[3] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[4]$_SDFFE_PN0P_  (.D(_00485_),
    .Q(\u_window_buffer.move_counter[4] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[5]$_SDFFE_PN0P_  (.D(_00486_),
    .Q(\u_window_buffer.move_counter[5] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[6]$_SDFFE_PN0P_  (.D(_00487_),
    .Q(\u_window_buffer.move_counter[6] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[7]$_SDFFE_PN0P_  (.D(_00488_),
    .Q(\u_window_buffer.move_counter[7] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[8]$_SDFFE_PN0P_  (.D(_00489_),
    .Q(\u_window_buffer.move_counter[8] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.move_counter[9]$_SDFFE_PN0P_  (.D(_00490_),
    .Q(\u_window_buffer.move_counter[9] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.next_state_is_valid_to_read$_DFF_P_  (.D(_00025_),
    .Q(\u_window_buffer.next_state_is_valid_to_read ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[0]$_SDFFE_PN0P_  (.D(_00491_),
    .Q(\u_window_buffer.read_ptr[0] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[10]$_SDFFE_PN0P_  (.D(_00492_),
    .Q(\u_window_buffer.read_ptr[10] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[11]$_SDFFE_PN0P_  (.D(_00493_),
    .Q(\u_window_buffer.read_ptr[11] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[12]$_SDFFE_PN0P_  (.D(_00494_),
    .Q(\u_window_buffer.read_ptr[12] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[13]$_SDFFE_PN0P_  (.D(_00495_),
    .Q(\u_window_buffer.read_ptr[13] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[14]$_SDFFE_PN0P_  (.D(_00496_),
    .Q(\u_window_buffer.read_ptr[14] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[15]$_SDFFE_PN0P_  (.D(_00497_),
    .Q(\u_window_buffer.read_ptr[15] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[16]$_SDFFE_PN0P_  (.D(_00498_),
    .Q(\u_window_buffer.read_ptr[16] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[17]$_SDFFE_PN0P_  (.D(_00499_),
    .Q(\u_window_buffer.read_ptr[17] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[18]$_SDFFE_PN0P_  (.D(_00500_),
    .Q(\u_window_buffer.read_ptr[18] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[19]$_SDFFE_PN0P_  (.D(_00501_),
    .Q(\u_window_buffer.read_ptr[19] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hs__dfxtp_4 \u_window_buffer.read_ptr[1]$_SDFFE_PN0P_  (.D(_00502_),
    .Q(\u_window_buffer.read_ptr[1] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[20]$_SDFFE_PN0P_  (.D(_00503_),
    .Q(\u_window_buffer.read_ptr[20] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[21]$_SDFFE_PN0P_  (.D(_00504_),
    .Q(\u_window_buffer.read_ptr[21] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[22]$_SDFFE_PN0P_  (.D(_00505_),
    .Q(\u_window_buffer.read_ptr[22] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[23]$_SDFFE_PN0P_  (.D(_00506_),
    .Q(\u_window_buffer.read_ptr[23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[24]$_SDFFE_PN0P_  (.D(_00507_),
    .Q(\u_window_buffer.read_ptr[24] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[25]$_SDFFE_PN0P_  (.D(_00508_),
    .Q(\u_window_buffer.read_ptr[25] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[26]$_SDFFE_PN0P_  (.D(_00509_),
    .Q(\u_window_buffer.read_ptr[26] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[27]$_SDFFE_PN0P_  (.D(_00510_),
    .Q(\u_window_buffer.read_ptr[27] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[28]$_SDFFE_PN0P_  (.D(_00511_),
    .Q(\u_window_buffer.read_ptr[28] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[29]$_SDFFE_PN0P_  (.D(_00512_),
    .Q(\u_window_buffer.read_ptr[29] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[2]$_SDFFE_PN0P_  (.D(_00513_),
    .Q(\u_window_buffer.read_ptr[2] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[30]$_SDFFE_PN0P_  (.D(_00514_),
    .Q(\u_window_buffer.read_ptr[30] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[31]$_SDFFE_PN0P_  (.D(_00515_),
    .Q(\u_window_buffer.read_ptr[31] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[3]$_SDFFE_PN0P_  (.D(_00516_),
    .Q(\u_window_buffer.read_ptr[3] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[4]$_SDFFE_PN0P_  (.D(_00517_),
    .Q(\u_window_buffer.read_ptr[4] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[5]$_SDFFE_PN0P_  (.D(_00518_),
    .Q(\u_window_buffer.read_ptr[5] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[6]$_SDFFE_PN0P_  (.D(_00519_),
    .Q(\u_window_buffer.read_ptr[6] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.read_ptr[7]$_SDFFE_PN0P_  (.D(_00520_),
    .Q(\u_window_buffer.read_ptr[7] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[8]$_SDFFE_PN0P_  (.D(_00521_),
    .Q(\u_window_buffer.read_ptr[8] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.read_ptr[9]$_SDFFE_PN0P_  (.D(_00522_),
    .Q(\u_window_buffer.read_ptr[9] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.start_next_state_o$_SDFF_PN0_  (.D(_00523_),
    .Q(start_hamming),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.write_ptr[0]$_SDFFE_PN0P_  (.D(_00524_),
    .Q(\u_window_buffer.write_ptr[0] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[10]$_SDFFE_PN0P_  (.D(_00525_),
    .Q(\u_window_buffer.write_ptr[10] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[11]$_SDFFE_PN0P_  (.D(_00526_),
    .Q(\u_window_buffer.write_ptr[11] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[12]$_SDFFE_PN0P_  (.D(_00527_),
    .Q(\u_window_buffer.write_ptr[12] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[13]$_SDFFE_PN0P_  (.D(_00528_),
    .Q(\u_window_buffer.write_ptr[13] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[14]$_SDFFE_PN0P_  (.D(_00529_),
    .Q(\u_window_buffer.write_ptr[14] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[15]$_SDFFE_PN0P_  (.D(_00530_),
    .Q(\u_window_buffer.write_ptr[15] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[16]$_SDFFE_PN0P_  (.D(_00531_),
    .Q(\u_window_buffer.write_ptr[16] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[17]$_SDFFE_PN0P_  (.D(_00532_),
    .Q(\u_window_buffer.write_ptr[17] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[18]$_SDFFE_PN0P_  (.D(_00533_),
    .Q(\u_window_buffer.write_ptr[18] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[19]$_SDFFE_PN0P_  (.D(_00534_),
    .Q(\u_window_buffer.write_ptr[19] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.write_ptr[1]$_SDFFE_PN0P_  (.D(_00535_),
    .Q(\u_window_buffer.write_ptr[1] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[20]$_SDFFE_PN0P_  (.D(_00536_),
    .Q(\u_window_buffer.write_ptr[20] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[21]$_SDFFE_PN0P_  (.D(_00537_),
    .Q(\u_window_buffer.write_ptr[21] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[22]$_SDFFE_PN0P_  (.D(_00538_),
    .Q(\u_window_buffer.write_ptr[22] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[23]$_SDFFE_PN0P_  (.D(_00539_),
    .Q(\u_window_buffer.write_ptr[23] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[24]$_SDFFE_PN0P_  (.D(_00540_),
    .Q(\u_window_buffer.write_ptr[24] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[25]$_SDFFE_PN0P_  (.D(_00541_),
    .Q(\u_window_buffer.write_ptr[25] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[26]$_SDFFE_PN0P_  (.D(_00542_),
    .Q(\u_window_buffer.write_ptr[26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[27]$_SDFFE_PN0P_  (.D(_00543_),
    .Q(\u_window_buffer.write_ptr[27] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[28]$_SDFFE_PN0P_  (.D(_00544_),
    .Q(\u_window_buffer.write_ptr[28] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[29]$_SDFFE_PN0P_  (.D(_00545_),
    .Q(\u_window_buffer.write_ptr[29] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hs__dfxtp_2 \u_window_buffer.write_ptr[2]$_SDFFE_PN0P_  (.D(_00546_),
    .Q(\u_window_buffer.write_ptr[2] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[30]$_SDFFE_PN0P_  (.D(_00547_),
    .Q(\u_window_buffer.write_ptr[30] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[31]$_SDFFE_PN0P_  (.D(_00548_),
    .Q(\u_window_buffer.write_ptr[31] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[3]$_SDFFE_PN0P_  (.D(_00549_),
    .Q(\u_window_buffer.write_ptr[3] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[4]$_SDFFE_PN0P_  (.D(_00550_),
    .Q(\u_window_buffer.write_ptr[4] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[5]$_SDFFE_PN0P_  (.D(_00551_),
    .Q(\u_window_buffer.write_ptr[5] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[6]$_SDFFE_PN0P_  (.D(_00552_),
    .Q(\u_window_buffer.write_ptr[6] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[7]$_SDFFE_PN0P_  (.D(_00553_),
    .Q(\u_window_buffer.write_ptr[7] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[8]$_SDFFE_PN0P_  (.D(_00554_),
    .Q(\u_window_buffer.write_ptr[8] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hs__dfxtp_1 \u_window_buffer.write_ptr[9]$_SDFFE_PN0P_  (.D(_00555_),
    .Q(\u_window_buffer.write_ptr[9] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hs__conb_1 _11643__1 (.LO(mfcc_data_o[0]));
 sky130_fd_sc_hs__conb_1 _11644__2 (.LO(mfcc_data_o[1]));
 sky130_fd_sc_hs__conb_1 _11645__3 (.LO(mfcc_data_o[2]));
 sky130_fd_sc_hs__conb_1 _11646__4 (.LO(mfcc_data_o[3]));
 sky130_fd_sc_hs__conb_1 _11647__5 (.LO(mfcc_data_o[4]));
 sky130_fd_sc_hs__conb_1 _11648__6 (.LO(mfcc_data_o[5]));
 sky130_fd_sc_hs__conb_1 _11649__7 (.LO(mfcc_data_o[6]));
 sky130_fd_sc_hs__conb_1 _11650__8 (.LO(mfcc_data_o[7]));
 sky130_fd_sc_hs__conb_1 _11651__9 (.LO(mfcc_data_o[8]));
 sky130_fd_sc_hs__conb_1 _11652__10 (.LO(mfcc_data_o[9]));
 sky130_fd_sc_hs__conb_1 _11653__11 (.LO(mfcc_data_o[10]));
 sky130_fd_sc_hs__conb_1 _11654__12 (.LO(mfcc_data_o[11]));
 sky130_fd_sc_hs__conb_1 _11655__13 (.LO(mfcc_data_o[12]));
 sky130_fd_sc_hs__conb_1 _11656__14 (.LO(mfcc_data_o[13]));
 sky130_fd_sc_hs__conb_1 _11657__15 (.LO(mfcc_data_o[14]));
 sky130_fd_sc_hs__conb_1 _11658__16 (.LO(mfcc_data_o[15]));
 sky130_fd_sc_hs__conb_1 _11659__17 (.LO(mfcc_data_o[16]));
 sky130_fd_sc_hs__conb_1 _11660__18 (.LO(mfcc_data_o[17]));
 sky130_fd_sc_hs__conb_1 _11661__19 (.LO(mfcc_data_o[18]));
 sky130_fd_sc_hs__conb_1 _11662__20 (.LO(mfcc_data_o[19]));
 sky130_fd_sc_hs__conb_1 _11663__21 (.LO(mfcc_data_o[20]));
 sky130_fd_sc_hs__conb_1 _11664__22 (.LO(mfcc_data_o[21]));
 sky130_fd_sc_hs__conb_1 _11665__23 (.LO(mfcc_data_o[22]));
 sky130_fd_sc_hs__conb_1 _11666__24 (.LO(mfcc_data_o[23]));
 sky130_fd_sc_hs__conb_1 _11667__25 (.LO(mfcc_data_o[24]));
 sky130_fd_sc_hs__conb_1 _11668__26 (.LO(mfcc_data_o[25]));
 sky130_fd_sc_hs__conb_1 _11669__27 (.LO(mfcc_data_o[26]));
 sky130_fd_sc_hs__conb_1 _11670__28 (.LO(mfcc_data_o[27]));
 sky130_fd_sc_hs__conb_1 _11671__29 (.LO(mfcc_data_o[28]));
 sky130_fd_sc_hs__conb_1 _11672__30 (.LO(mfcc_data_o[29]));
 sky130_fd_sc_hs__conb_1 _11673__31 (.LO(mfcc_data_o[30]));
 sky130_fd_sc_hs__conb_1 _11674__32 (.LO(mfcc_data_o[31]));
 sky130_fd_sc_hs__conb_1 _11675__33 (.LO(mfcc_data_o[32]));
 sky130_fd_sc_hs__conb_1 _11676__34 (.LO(mfcc_data_o[33]));
 sky130_fd_sc_hs__conb_1 _11677__35 (.LO(mfcc_data_o[34]));
 sky130_fd_sc_hs__conb_1 _11678__36 (.LO(mfcc_data_o[35]));
 sky130_fd_sc_hs__conb_1 _11679__37 (.LO(mfcc_data_o[36]));
 sky130_fd_sc_hs__conb_1 _11680__38 (.LO(mfcc_data_o[37]));
 sky130_fd_sc_hs__conb_1 _11681__39 (.LO(mfcc_data_o[38]));
 sky130_fd_sc_hs__conb_1 _11682__40 (.LO(mfcc_data_o[39]));
 sky130_fd_sc_hs__conb_1 _11683__41 (.LO(mfcc_data_o[40]));
 sky130_fd_sc_hs__conb_1 _11684__42 (.LO(mfcc_data_o[41]));
 sky130_fd_sc_hs__conb_1 _11685__43 (.LO(mfcc_data_o[42]));
 sky130_fd_sc_hs__conb_1 _11686__44 (.LO(mfcc_data_o[43]));
 sky130_fd_sc_hs__conb_1 _11687__45 (.LO(mfcc_data_o[44]));
 sky130_fd_sc_hs__conb_1 _11688__46 (.LO(mfcc_data_o[45]));
 sky130_fd_sc_hs__conb_1 _11689__47 (.LO(mfcc_data_o[46]));
 sky130_fd_sc_hs__conb_1 _11690__48 (.LO(mfcc_data_o[47]));
 sky130_fd_sc_hs__conb_1 _11691__49 (.LO(mfcc_data_o[48]));
 sky130_fd_sc_hs__conb_1 _11692__50 (.LO(mfcc_data_o[49]));
 sky130_fd_sc_hs__conb_1 _11693__51 (.LO(mfcc_data_o[50]));
 sky130_fd_sc_hs__conb_1 _11694__52 (.LO(mfcc_data_o[51]));
 sky130_fd_sc_hs__conb_1 _11695__53 (.LO(mfcc_data_o[52]));
 sky130_fd_sc_hs__conb_1 _11696__54 (.LO(mfcc_data_o[53]));
 sky130_fd_sc_hs__conb_1 _11697__55 (.LO(mfcc_data_o[54]));
 sky130_fd_sc_hs__conb_1 _11698__56 (.LO(mfcc_data_o[55]));
 sky130_fd_sc_hs__conb_1 _11699__57 (.LO(mfcc_data_o[56]));
 sky130_fd_sc_hs__conb_1 _11700__58 (.LO(mfcc_data_o[57]));
 sky130_fd_sc_hs__conb_1 _11701__59 (.LO(mfcc_data_o[58]));
 sky130_fd_sc_hs__conb_1 _11702__60 (.LO(mfcc_data_o[59]));
 sky130_fd_sc_hs__conb_1 _11703__61 (.LO(mfcc_data_o[60]));
 sky130_fd_sc_hs__conb_1 _11704__62 (.LO(mfcc_data_o[61]));
 sky130_fd_sc_hs__conb_1 _11705__63 (.LO(mfcc_data_o[62]));
 sky130_fd_sc_hs__conb_1 _11706__64 (.LO(mfcc_data_o[63]));
 sky130_fd_sc_hs__conb_1 _11707__65 (.LO(mfcc_data_o[64]));
 sky130_fd_sc_hs__conb_1 _11708__66 (.LO(mfcc_data_o[65]));
 sky130_fd_sc_hs__conb_1 _11709__67 (.LO(mfcc_data_o[66]));
 sky130_fd_sc_hs__conb_1 _11710__68 (.LO(mfcc_data_o[67]));
 sky130_fd_sc_hs__conb_1 _11711__69 (.LO(mfcc_data_o[68]));
 sky130_fd_sc_hs__conb_1 _11712__70 (.LO(mfcc_data_o[69]));
 sky130_fd_sc_hs__conb_1 _11713__71 (.LO(mfcc_data_o[70]));
 sky130_fd_sc_hs__conb_1 _11714__72 (.LO(mfcc_data_o[71]));
 sky130_fd_sc_hs__conb_1 _11715__73 (.LO(mfcc_data_o[72]));
 sky130_fd_sc_hs__conb_1 _11716__74 (.LO(mfcc_data_o[73]));
 sky130_fd_sc_hs__conb_1 _11717__75 (.LO(mfcc_data_o[74]));
 sky130_fd_sc_hs__conb_1 _11718__76 (.LO(mfcc_data_o[75]));
 sky130_fd_sc_hs__conb_1 _11719__77 (.LO(mfcc_data_o[76]));
 sky130_fd_sc_hs__conb_1 _11720__78 (.LO(mfcc_data_o[77]));
 sky130_fd_sc_hs__conb_1 _11721__79 (.LO(mfcc_data_o[78]));
 sky130_fd_sc_hs__conb_1 _11722__80 (.LO(mfcc_data_o[79]));
 sky130_fd_sc_hs__conb_1 _11723__81 (.LO(mfcc_data_o[80]));
 sky130_fd_sc_hs__conb_1 _11724__82 (.LO(mfcc_data_o[81]));
 sky130_fd_sc_hs__conb_1 _11725__83 (.LO(mfcc_data_o[82]));
 sky130_fd_sc_hs__conb_1 _11726__84 (.LO(mfcc_data_o[83]));
 sky130_fd_sc_hs__conb_1 _11727__85 (.LO(mfcc_data_o[84]));
 sky130_fd_sc_hs__conb_1 _11728__86 (.LO(mfcc_data_o[85]));
 sky130_fd_sc_hs__conb_1 _11729__87 (.LO(mfcc_data_o[86]));
 sky130_fd_sc_hs__conb_1 _11730__88 (.LO(mfcc_data_o[87]));
 sky130_fd_sc_hs__conb_1 _11731__89 (.LO(mfcc_data_o[88]));
 sky130_fd_sc_hs__conb_1 _11732__90 (.LO(mfcc_data_o[89]));
 sky130_fd_sc_hs__conb_1 _11733__91 (.LO(mfcc_data_o[90]));
 sky130_fd_sc_hs__conb_1 _11734__92 (.LO(mfcc_data_o[91]));
 sky130_fd_sc_hs__conb_1 _11735__93 (.LO(mfcc_data_o[92]));
 sky130_fd_sc_hs__conb_1 _11736__94 (.LO(mfcc_data_o[93]));
 sky130_fd_sc_hs__conb_1 _11737__95 (.LO(mfcc_data_o[94]));
 sky130_fd_sc_hs__conb_1 _11738__96 (.LO(mfcc_data_o[95]));
 sky130_fd_sc_hs__conb_1 _11739__97 (.LO(mfcc_data_o[96]));
 sky130_fd_sc_hs__conb_1 _11740__98 (.LO(mfcc_data_o[97]));
 sky130_fd_sc_hs__conb_1 _11741__99 (.LO(mfcc_data_o[98]));
 sky130_fd_sc_hs__conb_1 _11742__100 (.LO(mfcc_data_o[99]));
 sky130_fd_sc_hs__conb_1 _11743__101 (.LO(mfcc_data_o[100]));
 sky130_fd_sc_hs__conb_1 _11744__102 (.LO(mfcc_data_o[101]));
 sky130_fd_sc_hs__conb_1 _11745__103 (.LO(mfcc_data_o[102]));
 sky130_fd_sc_hs__conb_1 _11746__104 (.LO(mfcc_data_o[103]));
 sky130_fd_sc_hs__conb_1 _11747__105 (.LO(mfcc_data_o[104]));
 sky130_fd_sc_hs__conb_1 _11748__106 (.LO(mfcc_data_o[105]));
 sky130_fd_sc_hs__conb_1 _11749__107 (.LO(mfcc_data_o[106]));
 sky130_fd_sc_hs__conb_1 _11750__108 (.LO(mfcc_data_o[107]));
 sky130_fd_sc_hs__conb_1 _11751__109 (.LO(mfcc_data_o[108]));
 sky130_fd_sc_hs__conb_1 _11752__110 (.LO(mfcc_data_o[109]));
 sky130_fd_sc_hs__conb_1 _11753__111 (.LO(mfcc_data_o[110]));
 sky130_fd_sc_hs__conb_1 _11754__112 (.LO(mfcc_data_o[111]));
 sky130_fd_sc_hs__conb_1 _11755__113 (.LO(mfcc_data_o[112]));
 sky130_fd_sc_hs__conb_1 _11756__114 (.LO(mfcc_data_o[113]));
 sky130_fd_sc_hs__conb_1 _11757__115 (.LO(mfcc_data_o[114]));
 sky130_fd_sc_hs__conb_1 _11758__116 (.LO(mfcc_data_o[115]));
 sky130_fd_sc_hs__conb_1 _11759__117 (.LO(mfcc_data_o[116]));
 sky130_fd_sc_hs__conb_1 _11760__118 (.LO(mfcc_data_o[117]));
 sky130_fd_sc_hs__conb_1 _11761__119 (.LO(mfcc_data_o[118]));
 sky130_fd_sc_hs__conb_1 _11762__120 (.LO(mfcc_data_o[119]));
 sky130_fd_sc_hs__conb_1 _11763__121 (.LO(mfcc_data_o[120]));
 sky130_fd_sc_hs__conb_1 _11764__122 (.LO(mfcc_data_o[121]));
 sky130_fd_sc_hs__conb_1 _11765__123 (.LO(mfcc_data_o[122]));
 sky130_fd_sc_hs__conb_1 _11766__124 (.LO(mfcc_data_o[123]));
 sky130_fd_sc_hs__conb_1 _11767__125 (.LO(mfcc_data_o[124]));
 sky130_fd_sc_hs__conb_1 _11768__126 (.LO(mfcc_data_o[125]));
 sky130_fd_sc_hs__conb_1 _11769__127 (.LO(mfcc_data_o[126]));
 sky130_fd_sc_hs__conb_1 _11770__128 (.LO(mfcc_data_o[127]));
 sky130_fd_sc_hs__conb_1 _11771__129 (.LO(mfcc_data_o[128]));
 sky130_fd_sc_hs__conb_1 _11772__130 (.LO(mfcc_data_o[129]));
 sky130_fd_sc_hs__conb_1 _11773__131 (.LO(mfcc_data_o[130]));
 sky130_fd_sc_hs__conb_1 _11774__132 (.LO(mfcc_data_o[131]));
 sky130_fd_sc_hs__conb_1 _11775__133 (.LO(mfcc_data_o[132]));
 sky130_fd_sc_hs__conb_1 _11776__134 (.LO(mfcc_data_o[133]));
 sky130_fd_sc_hs__conb_1 _11777__135 (.LO(mfcc_data_o[134]));
 sky130_fd_sc_hs__conb_1 _11778__136 (.LO(mfcc_data_o[135]));
 sky130_fd_sc_hs__conb_1 _11779__137 (.LO(mfcc_data_o[136]));
 sky130_fd_sc_hs__conb_1 _11780__138 (.LO(mfcc_data_o[137]));
 sky130_fd_sc_hs__conb_1 _11781__139 (.LO(mfcc_data_o[138]));
 sky130_fd_sc_hs__conb_1 _11782__140 (.LO(mfcc_data_o[139]));
 sky130_fd_sc_hs__conb_1 _11783__141 (.LO(mfcc_data_o[140]));
 sky130_fd_sc_hs__conb_1 _11784__142 (.LO(mfcc_data_o[141]));
 sky130_fd_sc_hs__conb_1 _11785__143 (.LO(mfcc_data_o[142]));
 sky130_fd_sc_hs__conb_1 _11786__144 (.LO(mfcc_data_o[143]));
 sky130_fd_sc_hs__conb_1 _11787__145 (.LO(mfcc_data_o[144]));
 sky130_fd_sc_hs__conb_1 _11788__146 (.LO(mfcc_data_o[145]));
 sky130_fd_sc_hs__conb_1 _11789__147 (.LO(mfcc_data_o[146]));
 sky130_fd_sc_hs__conb_1 _11790__148 (.LO(mfcc_data_o[147]));
 sky130_fd_sc_hs__conb_1 _11791__149 (.LO(mfcc_data_o[148]));
 sky130_fd_sc_hs__conb_1 _11792__150 (.LO(mfcc_data_o[149]));
 sky130_fd_sc_hs__conb_1 _11793__151 (.LO(mfcc_data_o[150]));
 sky130_fd_sc_hs__conb_1 _11794__152 (.LO(mfcc_data_o[151]));
 sky130_fd_sc_hs__conb_1 _11795__153 (.LO(mfcc_data_o[152]));
 sky130_fd_sc_hs__conb_1 _11796__154 (.LO(mfcc_data_o[153]));
 sky130_fd_sc_hs__conb_1 _11797__155 (.LO(mfcc_data_o[154]));
 sky130_fd_sc_hs__conb_1 _11798__156 (.LO(mfcc_data_o[155]));
 sky130_fd_sc_hs__conb_1 _11799__157 (.LO(mfcc_data_o[156]));
 sky130_fd_sc_hs__conb_1 _11800__158 (.LO(mfcc_data_o[157]));
 sky130_fd_sc_hs__conb_1 _11801__159 (.LO(mfcc_data_o[158]));
 sky130_fd_sc_hs__conb_1 _11802__160 (.LO(mfcc_data_o[159]));
 sky130_fd_sc_hs__conb_1 _11803__161 (.LO(mfcc_data_o[160]));
 sky130_fd_sc_hs__conb_1 _11804__162 (.LO(mfcc_data_o[161]));
 sky130_fd_sc_hs__conb_1 _11805__163 (.LO(mfcc_data_o[162]));
 sky130_fd_sc_hs__conb_1 _11806__164 (.LO(mfcc_data_o[163]));
 sky130_fd_sc_hs__conb_1 _11807__165 (.LO(mfcc_data_o[164]));
 sky130_fd_sc_hs__conb_1 _11808__166 (.LO(mfcc_data_o[165]));
 sky130_fd_sc_hs__conb_1 _11809__167 (.LO(mfcc_data_o[166]));
 sky130_fd_sc_hs__conb_1 _11810__168 (.LO(mfcc_data_o[167]));
 sky130_fd_sc_hs__conb_1 _11811__169 (.LO(mfcc_data_o[168]));
 sky130_fd_sc_hs__conb_1 _11812__170 (.LO(mfcc_data_o[169]));
 sky130_fd_sc_hs__conb_1 _11813__171 (.LO(mfcc_data_o[170]));
 sky130_fd_sc_hs__conb_1 _11814__172 (.LO(mfcc_data_o[171]));
 sky130_fd_sc_hs__conb_1 _11815__173 (.LO(mfcc_data_o[172]));
 sky130_fd_sc_hs__conb_1 _11816__174 (.LO(mfcc_data_o[173]));
 sky130_fd_sc_hs__conb_1 _11817__175 (.LO(mfcc_data_o[174]));
 sky130_fd_sc_hs__conb_1 _11818__176 (.LO(mfcc_data_o[175]));
 sky130_fd_sc_hs__conb_1 _11819__177 (.LO(mfcc_data_o[176]));
 sky130_fd_sc_hs__conb_1 _11820__178 (.LO(mfcc_data_o[177]));
 sky130_fd_sc_hs__conb_1 _11821__179 (.LO(mfcc_data_o[178]));
 sky130_fd_sc_hs__conb_1 _11822__180 (.LO(mfcc_data_o[179]));
 sky130_fd_sc_hs__conb_1 _11823__181 (.LO(mfcc_data_o[180]));
 sky130_fd_sc_hs__conb_1 _11824__182 (.LO(mfcc_data_o[181]));
 sky130_fd_sc_hs__conb_1 _11825__183 (.LO(mfcc_data_o[182]));
 sky130_fd_sc_hs__conb_1 _11826__184 (.LO(mfcc_data_o[183]));
 sky130_fd_sc_hs__conb_1 _11827__185 (.LO(mfcc_data_o[184]));
 sky130_fd_sc_hs__conb_1 _11828__186 (.LO(mfcc_data_o[185]));
 sky130_fd_sc_hs__conb_1 _11829__187 (.LO(mfcc_data_o[186]));
 sky130_fd_sc_hs__conb_1 _11830__188 (.LO(mfcc_data_o[187]));
 sky130_fd_sc_hs__conb_1 _11831__189 (.LO(mfcc_data_o[188]));
 sky130_fd_sc_hs__conb_1 _11832__190 (.LO(mfcc_data_o[189]));
 sky130_fd_sc_hs__conb_1 _11833__191 (.LO(mfcc_data_o[190]));
 sky130_fd_sc_hs__conb_1 _11834__192 (.LO(mfcc_data_o[191]));
 sky130_fd_sc_hs__conb_1 _11835__193 (.LO(mfcc_data_o[192]));
 sky130_fd_sc_hs__conb_1 _11836__194 (.LO(mfcc_data_o[193]));
 sky130_fd_sc_hs__conb_1 _11837__195 (.LO(mfcc_data_o[194]));
 sky130_fd_sc_hs__conb_1 _11838__196 (.LO(mfcc_data_o[195]));
 sky130_fd_sc_hs__conb_1 _11839__197 (.LO(mfcc_data_o[196]));
 sky130_fd_sc_hs__conb_1 _11840__198 (.LO(mfcc_data_o[197]));
 sky130_fd_sc_hs__conb_1 _11841__199 (.LO(mfcc_data_o[198]));
 sky130_fd_sc_hs__conb_1 _11842__200 (.LO(mfcc_data_o[199]));
 sky130_fd_sc_hs__conb_1 _11843__201 (.LO(mfcc_data_o[200]));
 sky130_fd_sc_hs__conb_1 _11844__202 (.LO(mfcc_data_o[201]));
 sky130_fd_sc_hs__conb_1 _11845__203 (.LO(mfcc_data_o[202]));
 sky130_fd_sc_hs__conb_1 _11846__204 (.LO(mfcc_data_o[203]));
 sky130_fd_sc_hs__conb_1 _11847__205 (.LO(mfcc_data_o[204]));
 sky130_fd_sc_hs__conb_1 _11848__206 (.LO(mfcc_data_o[205]));
 sky130_fd_sc_hs__conb_1 _11849__207 (.LO(mfcc_data_o[206]));
 sky130_fd_sc_hs__conb_1 _11850__208 (.LO(mfcc_data_o[207]));
 sky130_fd_sc_hs__buf_1 rebuffer5096 (.A(_04842_),
    .X(net5096));
 sky130_fd_sc_hs__buf_1 place2198 (.A(_03457_),
    .X(net2198));
 sky130_fd_sc_hs__buf_1 place2200 (.A(_04540_),
    .X(net2200));
 sky130_fd_sc_hs__bufbuf_8 place2201 (.A(_04532_),
    .X(net2201));
 sky130_fd_sc_hs__buf_1 place2202 (.A(_04521_),
    .X(net2202));
 sky130_fd_sc_hs__buf_1 place2203 (.A(_04507_),
    .X(net2203));
 sky130_fd_sc_hs__buf_1 place2205 (.A(_01707_),
    .X(net2205));
 sky130_fd_sc_hs__buf_1 place2206 (.A(_01694_),
    .X(net2206));
 sky130_fd_sc_hs__buf_1 place2208 (.A(_05438_),
    .X(net2208));
 sky130_fd_sc_hs__clkbuf_2 place2209 (.A(_05419_),
    .X(net2209));
 sky130_fd_sc_hs__buf_1 place2210 (.A(_04530_),
    .X(net2210));
 sky130_fd_sc_hs__buf_1 place2211 (.A(_04499_),
    .X(net2211));
 sky130_fd_sc_hs__buf_1 place2212 (.A(_03458_),
    .X(net2212));
 sky130_fd_sc_hs__buf_1 place2213 (.A(_03431_),
    .X(net2213));
 sky130_fd_sc_hs__buf_1 place2215 (.A(_03414_),
    .X(net2215));
 sky130_fd_sc_hs__buf_1 place2216 (.A(_03401_),
    .X(net2216));
 sky130_fd_sc_hs__buf_1 place2217 (.A(_01675_),
    .X(net2217));
 sky130_fd_sc_hs__bufbuf_8 place2218 (.A(_01663_),
    .X(net2218));
 sky130_fd_sc_hs__buf_1 place2219 (.A(_05464_),
    .X(net2219));
 sky130_fd_sc_hs__bufbuf_8 place2220 (.A(_05424_),
    .X(net2220));
 sky130_fd_sc_hs__buf_1 place2221 (.A(_05410_),
    .X(net2221));
 sky130_fd_sc_hs__buf_1 place2222 (.A(_05400_),
    .X(net2222));
 sky130_fd_sc_hs__buf_1 place2224 (.A(_04500_),
    .X(net2224));
 sky130_fd_sc_hs__buf_1 place2226 (.A(_03399_),
    .X(net2226));
 sky130_fd_sc_hs__buf_1 place2225 (.A(_04498_),
    .X(net2225));
 sky130_fd_sc_hs__buf_1 place2227 (.A(_01677_),
    .X(net2227));
 sky130_fd_sc_hs__bufbuf_8 place2228 (.A(_05411_),
    .X(net2228));
 sky130_fd_sc_hs__buf_1 place2229 (.A(_05406_),
    .X(net2229));
 sky130_fd_sc_hs__buf_1 place2236 (.A(_03395_),
    .X(net2236));
 sky130_fd_sc_hs__buf_1 place2231 (.A(net5165),
    .X(net2231));
 sky130_fd_sc_hs__buf_1 place2232 (.A(_01657_),
    .X(net2232));
 sky130_fd_sc_hs__buf_1 place2233 (.A(_05399_),
    .X(net2233));
 sky130_fd_sc_hs__buf_1 place2234 (.A(_04494_),
    .X(net2234));
 sky130_fd_sc_hs__buf_1 place2235 (.A(_03398_),
    .X(net2235));
 sky130_fd_sc_hs__buf_1 place2238 (.A(_01656_),
    .X(net2238));
 sky130_fd_sc_hs__buf_1 place2240 (.A(_04505_),
    .X(net2240));
 sky130_fd_sc_hs__buf_1 place2242 (.A(_04486_),
    .X(net2242));
 sky130_fd_sc_hs__buf_1 place2243 (.A(_04478_),
    .X(net2243));
 sky130_fd_sc_hs__buf_2 place2245 (.A(_03400_),
    .X(net2245));
 sky130_fd_sc_hs__buf_1 place2246 (.A(_03394_),
    .X(net2246));
 sky130_fd_sc_hs__buf_1 place2247 (.A(_03389_),
    .X(net2247));
 sky130_fd_sc_hs__buf_1 place2248 (.A(_03378_),
    .X(net2248));
 sky130_fd_sc_hs__buf_1 place2251 (.A(_01649_),
    .X(net2251));
 sky130_fd_sc_hs__buf_1 place2249 (.A(_01665_),
    .X(net2249));
 sky130_fd_sc_hs__buf_1 place2250 (.A(_01664_),
    .X(net2250));
 sky130_fd_sc_hs__buf_1 place2252 (.A(_01641_),
    .X(net2252));
 sky130_fd_sc_hs__buf_1 place2253 (.A(_05397_),
    .X(net2253));
 sky130_fd_sc_hs__bufbuf_8 place2254 (.A(_04473_),
    .X(net2254));
 sky130_fd_sc_hs__buf_1 place2255 (.A(_03372_),
    .X(net2255));
 sky130_fd_sc_hs__buf_1 place2261 (.A(_05375_),
    .X(net2261));
 sky130_fd_sc_hs__buf_1 place2256 (.A(_01654_),
    .X(net2256));
 sky130_fd_sc_hs__buf_1 place2257 (.A(_01633_),
    .X(net2257));
 sky130_fd_sc_hs__buf_1 place2258 (.A(_05403_),
    .X(net2258));
 sky130_fd_sc_hs__buf_1 place2259 (.A(_05395_),
    .X(net2259));
 sky130_fd_sc_hs__buf_1 place2260 (.A(_05375_),
    .X(net2260));
 sky130_fd_sc_hs__buf_1 place2265 (.A(net2264),
    .X(net2265));
 sky130_fd_sc_hs__bufbuf_8 place2262 (.A(_04474_),
    .X(net2262));
 sky130_fd_sc_hs__buf_1 place2263 (.A(_04472_),
    .X(net2263));
 sky130_fd_sc_hs__buf_1 place2264 (.A(_03374_),
    .X(net2264));
 sky130_fd_sc_hs__buf_1 place2266 (.A(net4930),
    .X(net2266));
 sky130_fd_sc_hs__buf_1 place2268 (.A(_04469_),
    .X(net2268));
 sky130_fd_sc_hs__buf_1 place2267 (.A(_04469_),
    .X(net2267));
 sky130_fd_sc_hs__buf_1 place2269 (.A(_03390_),
    .X(net2269));
 sky130_fd_sc_hs__buf_1 place2270 (.A(net5139),
    .X(net2270));
 sky130_fd_sc_hs__buf_1 place2271 (.A(net5080),
    .X(net2271));
 sky130_fd_sc_hs__buf_1 place2272 (.A(_04471_),
    .X(net2272));
 sky130_fd_sc_hs__buf_1 place2274 (.A(_03392_),
    .X(net2274));
 sky130_fd_sc_hs__buf_1 place2277 (.A(_04459_),
    .X(net2277));
 sky130_fd_sc_hs__buf_1 place2278 (.A(_04451_),
    .X(net2278));
 sky130_fd_sc_hs__bufbuf_8 place2279 (.A(_03384_),
    .X(net2279));
 sky130_fd_sc_hs__buf_1 place2280 (.A(_03382_),
    .X(net2280));
 sky130_fd_sc_hs__buf_1 place2281 (.A(_03377_),
    .X(net2281));
 sky130_fd_sc_hs__buf_1 place2282 (.A(net5136),
    .X(net2282));
 sky130_fd_sc_hs__buf_1 place2283 (.A(_03357_),
    .X(net2283));
 sky130_fd_sc_hs__buf_1 place2284 (.A(_03348_),
    .X(net2284));
 sky130_fd_sc_hs__buf_1 place2285 (.A(_01621_),
    .X(net2285));
 sky130_fd_sc_hs__buf_1 place2286 (.A(_05380_),
    .X(net2286));
 sky130_fd_sc_hs__buf_2 place2287 (.A(_05353_),
    .X(net2287));
 sky130_fd_sc_hs__buf_2 place2289 (.A(_04463_),
    .X(net2289));
 sky130_fd_sc_hs__buf_1 place2290 (.A(_03369_),
    .X(net2290));
 sky130_fd_sc_hs__buf_1 place2291 (.A(_03343_),
    .X(net2291));
 sky130_fd_sc_hs__buf_1 place2292 (.A(_01639_),
    .X(net2292));
 sky130_fd_sc_hs__buf_1 place2293 (.A(_01606_),
    .X(net2293));
 sky130_fd_sc_hs__buf_1 place2296 (.A(net5072),
    .X(net2296));
 sky130_fd_sc_hs__buf_1 place2294 (.A(_05362_),
    .X(net2294));
 sky130_fd_sc_hs__buf_1 place2295 (.A(_05355_),
    .X(net2295));
 sky130_fd_sc_hs__buf_1 place2297 (.A(_04442_),
    .X(net2297));
 sky130_fd_sc_hs__buf_1 place2298 (.A(_03345_),
    .X(net2298));
 sky130_fd_sc_hs__buf_1 place2302 (.A(_05356_),
    .X(net2302));
 sky130_fd_sc_hs__buf_1 place2299 (.A(_01601_),
    .X(net2299));
 sky130_fd_sc_hs__buf_1 place2300 (.A(_01597_),
    .X(net2300));
 sky130_fd_sc_hs__buf_1 place2301 (.A(_05356_),
    .X(net2301));
 sky130_fd_sc_hs__buf_1 place2303 (.A(net4860),
    .X(net2303));
 sky130_fd_sc_hs__buf_1 place2304 (.A(net5177),
    .X(net2304));
 sky130_fd_sc_hs__buf_1 place2310 (.A(_03351_),
    .X(net2310));
 sky130_fd_sc_hs__buf_1 place2306 (.A(_01626_),
    .X(net2306));
 sky130_fd_sc_hs__buf_1 place2307 (.A(_01603_),
    .X(net2307));
 sky130_fd_sc_hs__bufbuf_8 place2309 (.A(_04467_),
    .X(net2309));
 sky130_fd_sc_hs__buf_1 place2308 (.A(_05339_),
    .X(net2308));
 sky130_fd_sc_hs__buf_1 place2311 (.A(_03322_),
    .X(net2311));
 sky130_fd_sc_hs__buf_1 place2312 (.A(_01611_),
    .X(net2312));
 sky130_fd_sc_hs__buf_1 place2315 (.A(_04446_),
    .X(net2315));
 sky130_fd_sc_hs__buf_1 place2317 (.A(_04430_),
    .X(net2317));
 sky130_fd_sc_hs__buf_1 place2318 (.A(_04421_),
    .X(net2318));
 sky130_fd_sc_hs__buf_1 place2319 (.A(_03338_),
    .X(net2319));
 sky130_fd_sc_hs__buf_1 place2320 (.A(net5196),
    .X(net2320));
 sky130_fd_sc_hs__buf_2 place2322 (.A(_01589_),
    .X(net2322));
 sky130_fd_sc_hs__buf_1 place2347 (.A(net2346),
    .X(net2347));
 sky130_fd_sc_hs__buf_1 place2323 (.A(net5101),
    .X(net2323));
 sky130_fd_sc_hs__buf_2 place2324 (.A(_05329_),
    .X(net2324));
 sky130_fd_sc_hs__buf_1 place2325 (.A(_05321_),
    .X(net2325));
 sky130_fd_sc_hs__buf_1 place2327 (.A(_04441_),
    .X(net2327));
 sky130_fd_sc_hs__buf_1 place2326 (.A(_04441_),
    .X(net2326));
 sky130_fd_sc_hs__buf_1 place2340 (.A(_04416_),
    .X(net2340));
 sky130_fd_sc_hs__buf_1 place2328 (.A(_04417_),
    .X(net2328));
 sky130_fd_sc_hs__buf_1 place2331 (.A(net2330),
    .X(net2331));
 sky130_fd_sc_hs__buf_4 place2329 (.A(_03341_),
    .X(net2329));
 sky130_fd_sc_hs__buf_1 place2330 (.A(_03332_),
    .X(net2330));
 sky130_fd_sc_hs__buf_1 place2339 (.A(_04416_),
    .X(net2339));
 sky130_fd_sc_hs__buf_1 place2332 (.A(_03321_),
    .X(net2332));
 sky130_fd_sc_hs__buf_1 place2335 (.A(net2334),
    .X(net2335));
 sky130_fd_sc_hs__buf_1 place2333 (.A(_01581_),
    .X(net2333));
 sky130_fd_sc_hs__buf_2 place2334 (.A(_05323_),
    .X(net2334));
 sky130_fd_sc_hs__buf_1 place2336 (.A(net5073),
    .X(net2336));
 sky130_fd_sc_hs__buf_1 place2337 (.A(_05306_),
    .X(net2337));
 sky130_fd_sc_hs__buf_1 place2338 (.A(_04418_),
    .X(net2338));
 sky130_fd_sc_hs__buf_1 place2345 (.A(_01566_),
    .X(net2345));
 sky130_fd_sc_hs__buf_1 place2341 (.A(_03331_),
    .X(net2341));
 sky130_fd_sc_hs__buf_1 place2342 (.A(_03323_),
    .X(net2342));
 sky130_fd_sc_hs__buf_1 place2343 (.A(_03315_),
    .X(net2343));
 sky130_fd_sc_hs__buf_1 place2344 (.A(_01594_),
    .X(net2344));
 sky130_fd_sc_hs__buf_1 place2346 (.A(_05325_),
    .X(net2346));
 sky130_fd_sc_hs__buf_1 place2348 (.A(_05313_),
    .X(net2348));
 sky130_fd_sc_hs__buf_1 place2351 (.A(net5175),
    .X(net2351));
 sky130_fd_sc_hs__buf_1 place2352 (.A(_01564_),
    .X(net2352));
 sky130_fd_sc_hs__buf_1 place2353 (.A(_05305_),
    .X(net2353));
 sky130_fd_sc_hs__buf_1 place2354 (.A(_04411_),
    .X(net2354));
 sky130_fd_sc_hs__buf_1 place2356 (.A(_03320_),
    .X(net2356));
 sky130_fd_sc_hs__buf_1 place2358 (.A(_05298_),
    .X(net2358));
 sky130_fd_sc_hs__buf_1 place2360 (.A(_04425_),
    .X(net2360));
 sky130_fd_sc_hs__buf_1 place2361 (.A(_04410_),
    .X(net2361));
 sky130_fd_sc_hs__buf_2 place2362 (.A(_04395_),
    .X(net2362));
 sky130_fd_sc_hs__buf_4 place2363 (.A(_03316_),
    .X(net2363));
 sky130_fd_sc_hs__buf_1 place2364 (.A(_03297_),
    .X(net2364));
 sky130_fd_sc_hs__buf_2 place2365 (.A(_03281_),
    .X(net2365));
 sky130_fd_sc_hs__buf_1 place2366 (.A(_01587_),
    .X(net2366));
 sky130_fd_sc_hs__buf_1 place2368 (.A(_01552_),
    .X(net2368));
 sky130_fd_sc_hs__buf_1 place2369 (.A(net4918),
    .X(net2369));
 sky130_fd_sc_hs__buf_1 place2370 (.A(_01537_),
    .X(net2370));
 sky130_fd_sc_hs__buf_1 place2371 (.A(_05342_),
    .X(net2371));
 sky130_fd_sc_hs__buf_1 place2375 (.A(_04401_),
    .X(net2375));
 sky130_fd_sc_hs__buf_1 place2376 (.A(_04391_),
    .X(net2376));
 sky130_fd_sc_hs__buf_1 place2384 (.A(net2383),
    .X(net2384));
 sky130_fd_sc_hs__buf_1 place2378 (.A(_03301_),
    .X(net2378));
 sky130_fd_sc_hs__buf_1 place2379 (.A(_03290_),
    .X(net2379));
 sky130_fd_sc_hs__buf_1 place2380 (.A(_03270_),
    .X(net2380));
 sky130_fd_sc_hs__buf_1 place2381 (.A(net4923),
    .X(net2381));
 sky130_fd_sc_hs__buf_2 place2382 (.A(_05302_),
    .X(net2382));
 sky130_fd_sc_hs__buf_1 place2383 (.A(_05279_),
    .X(net2383));
 sky130_fd_sc_hs__buf_1 place2387 (.A(_03298_),
    .X(net2387));
 sky130_fd_sc_hs__buf_1 place2385 (.A(_04402_),
    .X(net2385));
 sky130_fd_sc_hs__buf_1 place2386 (.A(_03300_),
    .X(net2386));
 sky130_fd_sc_hs__buf_1 place2388 (.A(_03277_),
    .X(net2388));
 sky130_fd_sc_hs__buf_1 place2390 (.A(_05286_),
    .X(net2390));
 sky130_fd_sc_hs__buf_1 place2389 (.A(_01525_),
    .X(net2389));
 sky130_fd_sc_hs__buf_1 place2391 (.A(_04381_),
    .X(net2391));
 sky130_fd_sc_hs__buf_1 place2393 (.A(_03309_),
    .X(net2393));
 sky130_fd_sc_hs__buf_1 place2396 (.A(_01548_),
    .X(net2396));
 sky130_fd_sc_hs__buf_1 rebuffer4923 (.A(_01547_),
    .X(net4923));
 sky130_fd_sc_hs__buf_1 place2398 (.A(_01523_),
    .X(net2398));
 sky130_fd_sc_hs__buf_1 place2397 (.A(_01523_),
    .X(net2397));
 sky130_fd_sc_hs__buf_1 place2401 (.A(_03280_),
    .X(net2401));
 sky130_fd_sc_hs__buf_1 place2399 (.A(net5082),
    .X(net2399));
 sky130_fd_sc_hs__buf_1 place2400 (.A(_04387_),
    .X(net2400));
 sky130_fd_sc_hs__buf_1 place2402 (.A(net5142),
    .X(net2402));
 sky130_fd_sc_hs__buf_2 place2403 (.A(net5181),
    .X(net2403));
 sky130_fd_sc_hs__buf_1 place2409 (.A(net2408),
    .X(net2409));
 sky130_fd_sc_hs__buf_1 place2404 (.A(_03255_),
    .X(net2404));
 sky130_fd_sc_hs__buf_1 place2405 (.A(net5192),
    .X(net2405));
 sky130_fd_sc_hs__buf_1 place2406 (.A(_01540_),
    .X(net2406));
 sky130_fd_sc_hs__buf_1 place2407 (.A(_01531_),
    .X(net2407));
 sky130_fd_sc_hs__buf_8 place2408 (.A(_01524_),
    .X(net2408));
 sky130_fd_sc_hs__buf_1 place2420 (.A(_01515_),
    .X(net2420));
 sky130_fd_sc_hs__bufbuf_8 place2412 (.A(_04379_),
    .X(net2412));
 sky130_fd_sc_hs__buf_1 place2410 (.A(net4919),
    .X(net2410));
 sky130_fd_sc_hs__buf_1 place2411 (.A(_04386_),
    .X(net2411));
 sky130_fd_sc_hs__buf_1 place2413 (.A(_04374_),
    .X(net2413));
 sky130_fd_sc_hs__buf_1 place2416 (.A(_03256_),
    .X(net2416));
 sky130_fd_sc_hs__buf_1 place2414 (.A(_04360_),
    .X(net2414));
 sky130_fd_sc_hs__buf_1 place2415 (.A(_03256_),
    .X(net2415));
 sky130_fd_sc_hs__buf_1 place2417 (.A(_01530_),
    .X(net2417));
 sky130_fd_sc_hs__buf_1 place2418 (.A(_01521_),
    .X(net2418));
 sky130_fd_sc_hs__buf_1 place2419 (.A(_01515_),
    .X(net2419));
 sky130_fd_sc_hs__buf_1 place2422 (.A(_01500_),
    .X(net2422));
 sky130_fd_sc_hs__buf_1 place2421 (.A(net4908),
    .X(net2421));
 sky130_fd_sc_hs__buf_2 place2423 (.A(_01496_),
    .X(net2423));
 sky130_fd_sc_hs__buf_1 place2424 (.A(_05283_),
    .X(net2424));
 sky130_fd_sc_hs__bufbuf_8 place2425 (.A(net5104),
    .X(net2425));
 sky130_fd_sc_hs__buf_1 place2426 (.A(_05269_),
    .X(net2426));
 sky130_fd_sc_hs__buf_1 place2427 (.A(_05262_),
    .X(net2427));
 sky130_fd_sc_hs__buf_1 place2429 (.A(_03262_),
    .X(net2429));
 sky130_fd_sc_hs__buf_1 place2430 (.A(_01499_),
    .X(net2430));
 sky130_fd_sc_hs__buf_1 place2444 (.A(_04351_),
    .X(net2444));
 sky130_fd_sc_hs__buf_2 place2433 (.A(net2432),
    .X(net2433));
 sky130_fd_sc_hs__buf_2 place2432 (.A(_05264_),
    .X(net2432));
 sky130_fd_sc_hs__buf_1 place2437 (.A(net2436),
    .X(net2437));
 sky130_fd_sc_hs__buf_1 place2434 (.A(_04354_),
    .X(net2434));
 sky130_fd_sc_hs__bufbuf_8 place2435 (.A(_03260_),
    .X(net2435));
 sky130_fd_sc_hs__buf_8 place2436 (.A(_03240_),
    .X(net2436));
 sky130_fd_sc_hs__bufbuf_8 place2438 (.A(_01503_),
    .X(net2438));
 sky130_fd_sc_hs__buf_1 place2439 (.A(_01492_),
    .X(net2439));
 sky130_fd_sc_hs__buf_1 place2442 (.A(_04375_),
    .X(net2442));
 sky130_fd_sc_hs__buf_2 place2440 (.A(_05266_),
    .X(net2440));
 sky130_fd_sc_hs__buf_1 place2441 (.A(_05251_),
    .X(net2441));
 sky130_fd_sc_hs__buf_1 place2443 (.A(_04353_),
    .X(net2443));
 sky130_fd_sc_hs__buf_1 place2445 (.A(_04341_),
    .X(net2445));
 sky130_fd_sc_hs__buf_1 place2447 (.A(_01483_),
    .X(net2447));
 sky130_fd_sc_hs__buf_1 place2448 (.A(_05247_),
    .X(net2448));
 sky130_fd_sc_hs__buf_1 place2450 (.A(_04364_),
    .X(net2450));
 sky130_fd_sc_hs__buf_1 place2451 (.A(_04350_),
    .X(net2451));
 sky130_fd_sc_hs__buf_1 place2501 (.A(_01477_),
    .X(net2501));
 sky130_fd_sc_hs__buf_1 place2453 (.A(_03261_),
    .X(net2453));
 sky130_fd_sc_hs__buf_1 place2454 (.A(_03251_),
    .X(net2454));
 sky130_fd_sc_hs__buf_1 place2455 (.A(_03250_),
    .X(net2455));
 sky130_fd_sc_hs__buf_1 place2456 (.A(_03237_),
    .X(net2456));
 sky130_fd_sc_hs__buf_1 place2457 (.A(net5172),
    .X(net2457));
 sky130_fd_sc_hs__buf_1 place2458 (.A(_03225_),
    .X(net2458));
 sky130_fd_sc_hs__buf_1 place2494 (.A(net2493),
    .X(net2494));
 sky130_fd_sc_hs__buf_1 place2459 (.A(_05222_),
    .X(net2459));
 sky130_fd_sc_hs__buf_1 place2483 (.A(net2482),
    .X(net2483));
 sky130_fd_sc_hs__buf_1 place2460 (.A(_04345_),
    .X(net2460));
 sky130_fd_sc_hs__bufbuf_8 place2461 (.A(_04342_),
    .X(net2461));
 sky130_fd_sc_hs__buf_1 place2462 (.A(_04335_),
    .X(net2462));
 sky130_fd_sc_hs__buf_1 place2463 (.A(_03232_),
    .X(net2463));
 sky130_fd_sc_hs__buf_2 place2464 (.A(_01495_),
    .X(net2464));
 sky130_fd_sc_hs__buf_1 place2468 (.A(_01462_),
    .X(net2468));
 sky130_fd_sc_hs__bufbuf_8 place2465 (.A(_01481_),
    .X(net2465));
 sky130_fd_sc_hs__buf_1 place2466 (.A(_01473_),
    .X(net2466));
 sky130_fd_sc_hs__buf_1 place2467 (.A(_01462_),
    .X(net2467));
 sky130_fd_sc_hs__buf_1 place2470 (.A(_05244_),
    .X(net2470));
 sky130_fd_sc_hs__buf_1 place2469 (.A(_05257_),
    .X(net2469));
 sky130_fd_sc_hs__buf_2 place2471 (.A(_05239_),
    .X(net2471));
 sky130_fd_sc_hs__buf_1 place2473 (.A(_04337_),
    .X(net2473));
 sky130_fd_sc_hs__buf_1 place2472 (.A(_05231_),
    .X(net2472));
 sky130_fd_sc_hs__buf_1 place2475 (.A(net2474),
    .X(net2475));
 sky130_fd_sc_hs__buf_4 place2474 (.A(_03241_),
    .X(net2474));
 sky130_fd_sc_hs__buf_2 place2480 (.A(_01456_),
    .X(net2480));
 sky130_fd_sc_hs__buf_1 place2476 (.A(_03234_),
    .X(net2476));
 sky130_fd_sc_hs__buf_1 rebuffer5142 (.A(_03275_),
    .X(net5142));
 sky130_fd_sc_hs__buf_1 place2477 (.A(_03224_),
    .X(net2477));
 sky130_fd_sc_hs__buf_1 place2479 (.A(_01456_),
    .X(net2479));
 sky130_fd_sc_hs__buf_2 place2482 (.A(_05225_),
    .X(net2482));
 sky130_fd_sc_hs__buf_1 place2481 (.A(_05225_),
    .X(net2481));
 sky130_fd_sc_hs__buf_1 place2484 (.A(_04330_),
    .X(net2484));
 sky130_fd_sc_hs__buf_1 place2491 (.A(_01451_),
    .X(net2491));
 sky130_fd_sc_hs__buf_1 place2485 (.A(net5115),
    .X(net2485));
 sky130_fd_sc_hs__buf_1 place2486 (.A(_01458_),
    .X(net2486));
 sky130_fd_sc_hs__buf_1 place2487 (.A(_01455_),
    .X(net2487));
 sky130_fd_sc_hs__buf_1 place2488 (.A(net5052),
    .X(net2488));
 sky130_fd_sc_hs__buf_1 place2489 (.A(_04339_),
    .X(net2489));
 sky130_fd_sc_hs__buf_1 place2490 (.A(_03212_),
    .X(net2490));
 sky130_fd_sc_hs__buf_1 place2492 (.A(net5045),
    .X(net2492));
 sky130_fd_sc_hs__buf_1 place2493 (.A(_04338_),
    .X(net2493));
 sky130_fd_sc_hs__buf_1 place2499 (.A(_03204_),
    .X(net2499));
 sky130_fd_sc_hs__bufbuf_8 place2495 (.A(_04328_),
    .X(net2495));
 sky130_fd_sc_hs__bufbuf_8 place2496 (.A(_04320_),
    .X(net2496));
 sky130_fd_sc_hs__buf_1 place2497 (.A(_03211_),
    .X(net2497));
 sky130_fd_sc_hs__buf_1 place2498 (.A(net5182),
    .X(net2498));
 sky130_fd_sc_hs__buf_1 place2500 (.A(_01506_),
    .X(net2500));
 sky130_fd_sc_hs__buf_1 place2503 (.A(_05210_),
    .X(net2503));
 sky130_fd_sc_hs__buf_2 place2507 (.A(_03189_),
    .X(net2507));
 sky130_fd_sc_hs__buf_1 place2509 (.A(_03183_),
    .X(net2509));
 sky130_fd_sc_hs__buf_1 place2510 (.A(_01461_),
    .X(net2510));
 sky130_fd_sc_hs__buf_1 place2511 (.A(_01449_),
    .X(net2511));
 sky130_fd_sc_hs__buf_1 place2512 (.A(_01432_),
    .X(net2512));
 sky130_fd_sc_hs__buf_1 place2513 (.A(_05234_),
    .X(net2513));
 sky130_fd_sc_hs__buf_1 place2515 (.A(_05201_),
    .X(net2515));
 sky130_fd_sc_hs__buf_1 place2516 (.A(_05193_),
    .X(net2516));
 sky130_fd_sc_hs__buf_1 place2518 (.A(_03193_),
    .X(net2518));
 sky130_fd_sc_hs__buf_1 place2519 (.A(_01454_),
    .X(net2519));
 sky130_fd_sc_hs__bufbuf_8 place2520 (.A(_01437_),
    .X(net2520));
 sky130_fd_sc_hs__buf_1 place2522 (.A(_05215_),
    .X(net2522));
 sky130_fd_sc_hs__buf_1 place2521 (.A(_05215_),
    .X(net2521));
 sky130_fd_sc_hs__buf_1 place2523 (.A(_05188_),
    .X(net2523));
 sky130_fd_sc_hs__buf_1 place2525 (.A(_04299_),
    .X(net2525));
 sky130_fd_sc_hs__buf_2 place2524 (.A(_04299_),
    .X(net2524));
 sky130_fd_sc_hs__buf_1 place2536 (.A(_05184_),
    .X(net2536));
 sky130_fd_sc_hs__buf_1 place2526 (.A(net5113),
    .X(net2526));
 sky130_fd_sc_hs__buf_1 place2527 (.A(_01427_),
    .X(net2527));
 sky130_fd_sc_hs__buf_8 clone4961 (.A(_04787_),
    .X(net4961));
 sky130_fd_sc_hs__buf_1 place2535 (.A(_05184_),
    .X(net2535));
 sky130_fd_sc_hs__buf_1 place2529 (.A(_05189_),
    .X(net2529));
 sky130_fd_sc_hs__buf_1 place2530 (.A(_05187_),
    .X(net2530));
 sky130_fd_sc_hs__buf_1 place2531 (.A(_04321_),
    .X(net2531));
 sky130_fd_sc_hs__buf_1 place2532 (.A(_03210_),
    .X(net2532));
 sky130_fd_sc_hs__buf_1 place2533 (.A(_01418_),
    .X(net2533));
 sky130_fd_sc_hs__buf_1 place2534 (.A(_05205_),
    .X(net2534));
 sky130_fd_sc_hs__buf_1 place2542 (.A(_03185_),
    .X(net2542));
 sky130_fd_sc_hs__buf_1 place2538 (.A(_04297_),
    .X(net2538));
 sky130_fd_sc_hs__buf_1 place2539 (.A(_04292_),
    .X(net2539));
 sky130_fd_sc_hs__buf_1 place2540 (.A(_04280_),
    .X(net2540));
 sky130_fd_sc_hs__buf_1 place2541 (.A(_03186_),
    .X(net2541));
 sky130_fd_sc_hs__buf_1 place2543 (.A(net5179),
    .X(net2543));
 sky130_fd_sc_hs__buf_1 place2544 (.A(_01431_),
    .X(net2544));
 sky130_fd_sc_hs__buf_1 place2546 (.A(_05204_),
    .X(net2546));
 sky130_fd_sc_hs__buf_2 place2547 (.A(_04273_),
    .X(net2547));
 sky130_fd_sc_hs__buf_1 place2556 (.A(net2555),
    .X(net2556));
 sky130_fd_sc_hs__buf_1 place2550 (.A(_03160_),
    .X(net2550));
 sky130_fd_sc_hs__buf_1 place2548 (.A(_03171_),
    .X(net2548));
 sky130_fd_sc_hs__buf_1 place2549 (.A(_03160_),
    .X(net2549));
 sky130_fd_sc_hs__buf_1 place2551 (.A(_01430_),
    .X(net2551));
 sky130_fd_sc_hs__buf_1 place2552 (.A(_01416_),
    .X(net2552));
 sky130_fd_sc_hs__buf_1 place2553 (.A(_01399_),
    .X(net2553));
 sky130_fd_sc_hs__buf_1 place2554 (.A(_05191_),
    .X(net2554));
 sky130_fd_sc_hs__buf_2 place2555 (.A(_05182_),
    .X(net2555));
 sky130_fd_sc_hs__buf_1 place2557 (.A(_05166_),
    .X(net2557));
 sky130_fd_sc_hs__buf_1 place2578 (.A(_05170_),
    .X(net2578));
 sky130_fd_sc_hs__buf_2 place2558 (.A(_04275_),
    .X(net2558));
 sky130_fd_sc_hs__buf_1 place2577 (.A(_01387_),
    .X(net2577));
 sky130_fd_sc_hs__clkbuf_2 place2565 (.A(_05159_),
    .X(net2565));
 sky130_fd_sc_hs__buf_1 place2559 (.A(_04272_),
    .X(net2559));
 sky130_fd_sc_hs__buf_1 place2560 (.A(_03179_),
    .X(net2560));
 sky130_fd_sc_hs__buf_2 place2561 (.A(_03173_),
    .X(net2561));
 sky130_fd_sc_hs__buf_1 place2562 (.A(_01405_),
    .X(net2562));
 sky130_fd_sc_hs__buf_1 place2563 (.A(_01392_),
    .X(net2563));
 sky130_fd_sc_hs__buf_1 place2564 (.A(_05186_),
    .X(net2564));
 sky130_fd_sc_hs__buf_1 place2570 (.A(net5047),
    .X(net2570));
 sky130_fd_sc_hs__buf_1 place2566 (.A(_04268_),
    .X(net2566));
 sky130_fd_sc_hs__buf_1 place2567 (.A(_01423_),
    .X(net2567));
 sky130_fd_sc_hs__buf_1 place2568 (.A(_01394_),
    .X(net2568));
 sky130_fd_sc_hs__buf_1 place2569 (.A(_01391_),
    .X(net2569));
 sky130_fd_sc_hs__buf_1 place2571 (.A(_05160_),
    .X(net2571));
 sky130_fd_sc_hs__buf_1 place2576 (.A(_03144_),
    .X(net2576));
 sky130_fd_sc_hs__buf_1 place2572 (.A(_05158_),
    .X(net2572));
 sky130_fd_sc_hs__buf_1 place2573 (.A(_04281_),
    .X(net2573));
 sky130_fd_sc_hs__bufbuf_8 place2574 (.A(_04279_),
    .X(net2574));
 sky130_fd_sc_hs__buf_1 place2575 (.A(_04267_),
    .X(net2575));
 sky130_fd_sc_hs__buf_1 place2579 (.A(net5079),
    .X(net2579));
 sky130_fd_sc_hs__buf_1 place2580 (.A(net5067),
    .X(net2580));
 sky130_fd_sc_hs__buf_1 place2581 (.A(_04285_),
    .X(net2581));
 sky130_fd_sc_hs__buf_1 place2583 (.A(_04271_),
    .X(net2583));
 sky130_fd_sc_hs__buf_1 place2584 (.A(_04259_),
    .X(net2584));
 sky130_fd_sc_hs__buf_1 place2585 (.A(_04248_),
    .X(net2585));
 sky130_fd_sc_hs__buf_1 place2586 (.A(_03194_),
    .X(net2586));
 sky130_fd_sc_hs__buf_1 place2587 (.A(_03150_),
    .X(net2587));
 sky130_fd_sc_hs__buf_1 place2588 (.A(_01420_),
    .X(net2588));
 sky130_fd_sc_hs__buf_1 place2590 (.A(_04270_),
    .X(net2590));
 sky130_fd_sc_hs__buf_1 place2589 (.A(_05174_),
    .X(net2589));
 sky130_fd_sc_hs__buf_1 place2634 (.A(_01364_),
    .X(net2634));
 sky130_fd_sc_hs__buf_1 place2592 (.A(_03156_),
    .X(net2592));
 sky130_fd_sc_hs__buf_1 place2593 (.A(_03147_),
    .X(net2593));
 sky130_fd_sc_hs__buf_1 place2613 (.A(_01360_),
    .X(net2613));
 sky130_fd_sc_hs__bufbuf_8 place2594 (.A(_01419_),
    .X(net2594));
 sky130_fd_sc_hs__buf_2 place2595 (.A(_01398_),
    .X(net2595));
 sky130_fd_sc_hs__buf_1 place2596 (.A(_01390_),
    .X(net2596));
 sky130_fd_sc_hs__bufbuf_8 place2609 (.A(net5048),
    .X(net2609));
 sky130_fd_sc_hs__buf_1 place2599 (.A(_01367_),
    .X(net2599));
 sky130_fd_sc_hs__buf_2 place2597 (.A(_01385_),
    .X(net2597));
 sky130_fd_sc_hs__buf_1 place2598 (.A(_01367_),
    .X(net2598));
 sky130_fd_sc_hs__buf_1 place2600 (.A(_05164_),
    .X(net2600));
 sky130_fd_sc_hs__buf_1 place2606 (.A(net4863),
    .X(net2606));
 sky130_fd_sc_hs__buf_1 place2605 (.A(_01389_),
    .X(net2605));
 sky130_fd_sc_hs__buf_2 place2601 (.A(_05136_),
    .X(net2601));
 sky130_fd_sc_hs__buf_1 place2602 (.A(_04243_),
    .X(net2602));
 sky130_fd_sc_hs__buf_1 place2603 (.A(_03139_),
    .X(net2603));
 sky130_fd_sc_hs__buf_1 place2604 (.A(_01389_),
    .X(net2604));
 sky130_fd_sc_hs__buf_1 place2607 (.A(_01361_),
    .X(net2607));
 sky130_fd_sc_hs__buf_1 place2608 (.A(_05156_),
    .X(net2608));
 sky130_fd_sc_hs__buf_1 place2610 (.A(_05129_),
    .X(net2610));
 sky130_fd_sc_hs__buf_1 place2611 (.A(_04239_),
    .X(net2611));
 sky130_fd_sc_hs__buf_1 place2612 (.A(_03130_),
    .X(net2612));
 sky130_fd_sc_hs__buf_1 place2614 (.A(_04251_),
    .X(net2614));
 sky130_fd_sc_hs__buf_1 place2615 (.A(_04231_),
    .X(net2615));
 sky130_fd_sc_hs__buf_1 place2616 (.A(_01366_),
    .X(net2616));
 sky130_fd_sc_hs__buf_1 place2633 (.A(_01364_),
    .X(net2633));
 sky130_fd_sc_hs__buf_1 place2617 (.A(_05124_),
    .X(net2617));
 sky130_fd_sc_hs__bufbuf_8 place2618 (.A(_04252_),
    .X(net2618));
 sky130_fd_sc_hs__buf_1 place2619 (.A(_04247_),
    .X(net2619));
 sky130_fd_sc_hs__buf_1 place2631 (.A(_03096_),
    .X(net2631));
 sky130_fd_sc_hs__buf_1 place2620 (.A(_04238_),
    .X(net2620));
 sky130_fd_sc_hs__buf_1 place2621 (.A(_04230_),
    .X(net2621));
 sky130_fd_sc_hs__buf_1 place2622 (.A(_04221_),
    .X(net2622));
 sky130_fd_sc_hs__buf_1 place2623 (.A(_03136_),
    .X(net2623));
 sky130_fd_sc_hs__buf_1 place2630 (.A(_03114_),
    .X(net2630));
 sky130_fd_sc_hs__buf_1 place2624 (.A(net5141),
    .X(net2624));
 sky130_fd_sc_hs__buf_1 place2625 (.A(_03104_),
    .X(net2625));
 sky130_fd_sc_hs__buf_4 place2627 (.A(_04242_),
    .X(net2627));
 sky130_fd_sc_hs__buf_1 place2626 (.A(_05131_),
    .X(net2626));
 sky130_fd_sc_hs__buf_1 place2628 (.A(_04232_),
    .X(net2628));
 sky130_fd_sc_hs__buf_1 place2629 (.A(_04219_),
    .X(net2629));
 sky130_fd_sc_hs__buf_1 place2632 (.A(_01364_),
    .X(net2632));
 sky130_fd_sc_hs__buf_1 place2635 (.A(net4897),
    .X(net2635));
 sky130_fd_sc_hs__buf_1 place2637 (.A(_05146_),
    .X(net2637));
 sky130_fd_sc_hs__buf_1 place2636 (.A(_01335_),
    .X(net2636));
 sky130_fd_sc_hs__buf_1 place2638 (.A(_05115_),
    .X(net2638));
 sky130_fd_sc_hs__buf_2 place2644 (.A(_05120_),
    .X(net2644));
 sky130_fd_sc_hs__buf_1 place2640 (.A(_04233_),
    .X(net2640));
 sky130_fd_sc_hs__buf_1 place2641 (.A(_03115_),
    .X(net2641));
 sky130_fd_sc_hs__buf_1 place2642 (.A(net5143),
    .X(net2642));
 sky130_fd_sc_hs__buf_2 place2643 (.A(_01329_),
    .X(net2643));
 sky130_fd_sc_hs__buf_1 place2647 (.A(_04213_),
    .X(net2647));
 sky130_fd_sc_hs__bufbuf_8 place2645 (.A(_04226_),
    .X(net2645));
 sky130_fd_sc_hs__buf_1 place2646 (.A(_04213_),
    .X(net2646));
 sky130_fd_sc_hs__buf_1 place2649 (.A(_01358_),
    .X(net2649));
 sky130_fd_sc_hs__buf_1 place2648 (.A(_03095_),
    .X(net2648));
 sky130_fd_sc_hs__buf_1 place2651 (.A(_01331_),
    .X(net2651));
 sky130_fd_sc_hs__buf_1 place2652 (.A(_01328_),
    .X(net2652));
 sky130_fd_sc_hs__buf_1 place2653 (.A(_05137_),
    .X(net2653));
 sky130_fd_sc_hs__buf_1 place2656 (.A(net5097),
    .X(net2656));
 sky130_fd_sc_hs__buf_1 place2664 (.A(_04191_),
    .X(net2664));
 sky130_fd_sc_hs__bufbuf_8 place2657 (.A(_04225_),
    .X(net2657));
 sky130_fd_sc_hs__buf_2 place2658 (.A(_04212_),
    .X(net2658));
 sky130_fd_sc_hs__buf_1 place2659 (.A(_04197_),
    .X(net2659));
 sky130_fd_sc_hs__bufbuf_8 place2660 (.A(_03108_),
    .X(net2660));
 sky130_fd_sc_hs__buf_1 place2661 (.A(net5066),
    .X(net2661));
 sky130_fd_sc_hs__buf_1 place2662 (.A(_04203_),
    .X(net2662));
 sky130_fd_sc_hs__buf_1 place2663 (.A(_04191_),
    .X(net2663));
 sky130_fd_sc_hs__buf_1 place2666 (.A(_03092_),
    .X(net2666));
 sky130_fd_sc_hs__buf_1 place2667 (.A(_03083_),
    .X(net2667));
 sky130_fd_sc_hs__buf_1 place2669 (.A(_03075_),
    .X(net2669));
 sky130_fd_sc_hs__buf_1 place2675 (.A(_03065_),
    .X(net2675));
 sky130_fd_sc_hs__buf_1 place2674 (.A(_03065_),
    .X(net2674));
 sky130_fd_sc_hs__buf_1 place2671 (.A(_04192_),
    .X(net2671));
 sky130_fd_sc_hs__buf_1 place2670 (.A(_05089_),
    .X(net2670));
 sky130_fd_sc_hs__buf_1 place2672 (.A(_04190_),
    .X(net2672));
 sky130_fd_sc_hs__buf_1 place2673 (.A(_03067_),
    .X(net2673));
 sky130_fd_sc_hs__buf_2 place2676 (.A(_01374_),
    .X(net2676));
 sky130_fd_sc_hs__buf_1 place2678 (.A(_01334_),
    .X(net2678));
 sky130_fd_sc_hs__buf_1 place2679 (.A(_01322_),
    .X(net2679));
 sky130_fd_sc_hs__buf_1 place2681 (.A(net4907),
    .X(net2681));
 sky130_fd_sc_hs__bufbuf_8 place2682 (.A(_05111_),
    .X(net2682));
 sky130_fd_sc_hs__buf_1 place2683 (.A(_05095_),
    .X(net2683));
 sky130_fd_sc_hs__buf_1 place2686 (.A(_05080_),
    .X(net2686));
 sky130_fd_sc_hs__buf_1 place2687 (.A(_04186_),
    .X(net2687));
 sky130_fd_sc_hs__buf_1 place2688 (.A(_03066_),
    .X(net2688));
 sky130_fd_sc_hs__buf_1 place2689 (.A(_01337_),
    .X(net2689));
 sky130_fd_sc_hs__buf_1 place2691 (.A(_01299_),
    .X(net2691));
 sky130_fd_sc_hs__buf_2 place2692 (.A(_05090_),
    .X(net2692));
 sky130_fd_sc_hs__buf_1 place2695 (.A(net5116),
    .X(net2695));
 sky130_fd_sc_hs__buf_1 place2696 (.A(_01336_),
    .X(net2696));
 sky130_fd_sc_hs__buf_1 place2697 (.A(net4924),
    .X(net2697));
 sky130_fd_sc_hs__buf_1 place2698 (.A(_01301_),
    .X(net2698));
 sky130_fd_sc_hs__buf_1 place2712 (.A(_04189_),
    .X(net2712));
 sky130_fd_sc_hs__buf_1 place2699 (.A(_01298_),
    .X(net2699));
 sky130_fd_sc_hs__buf_1 place2700 (.A(_05098_),
    .X(net2700));
 sky130_fd_sc_hs__buf_1 place2701 (.A(_05091_),
    .X(net2701));
 sky130_fd_sc_hs__buf_1 place2708 (.A(_01297_),
    .X(net2708));
 sky130_fd_sc_hs__buf_1 place2702 (.A(_05079_),
    .X(net2702));
 sky130_fd_sc_hs__buf_1 place2703 (.A(_04195_),
    .X(net2703));
 sky130_fd_sc_hs__buf_1 place2704 (.A(_04178_),
    .X(net2704));
 sky130_fd_sc_hs__buf_1 place2705 (.A(_04169_),
    .X(net2705));
 sky130_fd_sc_hs__bufbuf_8 place2706 (.A(_03079_),
    .X(net2706));
 sky130_fd_sc_hs__buf_1 place2707 (.A(_03041_),
    .X(net2707));
 sky130_fd_sc_hs__buf_1 place2709 (.A(_01290_),
    .X(net2709));
 sky130_fd_sc_hs__buf_1 place2710 (.A(_05073_),
    .X(net2710));
 sky130_fd_sc_hs__buf_1 place2711 (.A(_04189_),
    .X(net2711));
 sky130_fd_sc_hs__buf_1 place2713 (.A(_04184_),
    .X(net2713));
 sky130_fd_sc_hs__buf_1 place2714 (.A(_04163_),
    .X(net2714));
 sky130_fd_sc_hs__buf_1 place2715 (.A(_03073_),
    .X(net2715));
 sky130_fd_sc_hs__buf_1 place2716 (.A(_03061_),
    .X(net2716));
 sky130_fd_sc_hs__buf_2 place2717 (.A(_03055_),
    .X(net2717));
 sky130_fd_sc_hs__buf_1 place2718 (.A(_03048_),
    .X(net2718));
 sky130_fd_sc_hs__bufbuf_8 place2719 (.A(_01316_),
    .X(net2719));
 sky130_fd_sc_hs__buf_1 place2720 (.A(_01315_),
    .X(net2720));
 sky130_fd_sc_hs__buf_1 place2721 (.A(_05082_),
    .X(net2721));
 sky130_fd_sc_hs__buf_1 place2723 (.A(_04164_),
    .X(net2723));
 sky130_fd_sc_hs__buf_1 place2724 (.A(_04162_),
    .X(net2724));
 sky130_fd_sc_hs__bufbuf_8 place2725 (.A(_01304_),
    .X(net2725));
 sky130_fd_sc_hs__buf_4 place2726 (.A(_01289_),
    .X(net2726));
 sky130_fd_sc_hs__buf_1 place2727 (.A(_01274_),
    .X(net2727));
 sky130_fd_sc_hs__buf_1 place2728 (.A(_05081_),
    .X(net2728));
 sky130_fd_sc_hs__buf_1 place2729 (.A(_05072_),
    .X(net2729));
 sky130_fd_sc_hs__buf_1 place2731 (.A(_04157_),
    .X(net2731));
 sky130_fd_sc_hs__buf_1 place2732 (.A(_03035_),
    .X(net2732));
 sky130_fd_sc_hs__buf_1 place2733 (.A(_05076_),
    .X(net2733));
 sky130_fd_sc_hs__buf_1 place2735 (.A(_05066_),
    .X(net2735));
 sky130_fd_sc_hs__buf_1 place2736 (.A(_05042_),
    .X(net2736));
 sky130_fd_sc_hs__buf_1 place2738 (.A(net5125),
    .X(net2738));
 sky130_fd_sc_hs__buf_1 place2739 (.A(_01282_),
    .X(net2739));
 sky130_fd_sc_hs__buf_1 place2743 (.A(_04204_),
    .X(net2743));
 sky130_fd_sc_hs__buf_1 place2740 (.A(_05064_),
    .X(net2740));
 sky130_fd_sc_hs__buf_1 place2741 (.A(_05044_),
    .X(net2741));
 sky130_fd_sc_hs__buf_1 place2742 (.A(net5053),
    .X(net2742));
 sky130_fd_sc_hs__buf_1 place2744 (.A(_04168_),
    .X(net2744));
 sky130_fd_sc_hs__buf_1 place2745 (.A(_04155_),
    .X(net2745));
 sky130_fd_sc_hs__buf_2 place2746 (.A(_04138_),
    .X(net2746));
 sky130_fd_sc_hs__buf_1 place2747 (.A(_03037_),
    .X(net2747));
 sky130_fd_sc_hs__buf_1 place2748 (.A(_03030_),
    .X(net2748));
 sky130_fd_sc_hs__bufbuf_8 place2750 (.A(_04145_),
    .X(net2750));
 sky130_fd_sc_hs__buf_1 place2751 (.A(_04129_),
    .X(net2751));
 sky130_fd_sc_hs__bufbuf_8 place2752 (.A(_03036_),
    .X(net2752));
 sky130_fd_sc_hs__buf_1 place2753 (.A(net5194),
    .X(net2753));
 sky130_fd_sc_hs__buf_1 place2755 (.A(net5169),
    .X(net2755));
 sky130_fd_sc_hs__buf_1 place2756 (.A(net5132),
    .X(net2756));
 sky130_fd_sc_hs__buf_1 place2757 (.A(net5069),
    .X(net2757));
 sky130_fd_sc_hs__buf_1 place2758 (.A(_04130_),
    .X(net2758));
 sky130_fd_sc_hs__buf_1 place2760 (.A(_03009_),
    .X(net2760));
 sky130_fd_sc_hs__buf_4 place2763 (.A(_01259_),
    .X(net2763));
 sky130_fd_sc_hs__buf_1 place2765 (.A(_01238_),
    .X(net2765));
 sky130_fd_sc_hs__bufbuf_8 place2766 (.A(_05049_),
    .X(net2766));
 sky130_fd_sc_hs__buf_1 place2767 (.A(net5092),
    .X(net2767));
 sky130_fd_sc_hs__buf_1 place2768 (.A(_04141_),
    .X(net2768));
 sky130_fd_sc_hs__buf_1 place2770 (.A(_03011_),
    .X(net2770));
 sky130_fd_sc_hs__buf_1 place2772 (.A(_01263_),
    .X(net2772));
 sky130_fd_sc_hs__buf_1 place2773 (.A(_01248_),
    .X(net2773));
 sky130_fd_sc_hs__buf_1 place2774 (.A(_01231_),
    .X(net2774));
 sky130_fd_sc_hs__buf_2 place2782 (.A(_05040_),
    .X(net2782));
 sky130_fd_sc_hs__buf_1 place2784 (.A(_05030_),
    .X(net2784));
 sky130_fd_sc_hs__buf_2 place2785 (.A(_05028_),
    .X(net2785));
 sky130_fd_sc_hs__buf_1 place2787 (.A(_04114_),
    .X(net2787));
 sky130_fd_sc_hs__bufbuf_8 place2789 (.A(_03023_),
    .X(net2789));
 sky130_fd_sc_hs__buf_1 place2790 (.A(_03016_),
    .X(net2790));
 sky130_fd_sc_hs__buf_1 place2791 (.A(_02996_),
    .X(net2791));
 sky130_fd_sc_hs__buf_2 place2797 (.A(_03002_),
    .X(net2797));
 sky130_fd_sc_hs__buf_1 place2793 (.A(_05012_),
    .X(net2793));
 sky130_fd_sc_hs__buf_1 place2794 (.A(_04123_),
    .X(net2794));
 sky130_fd_sc_hs__buf_1 place2795 (.A(_03015_),
    .X(net2795));
 sky130_fd_sc_hs__buf_1 place2796 (.A(_03007_),
    .X(net2796));
 sky130_fd_sc_hs__buf_1 place2798 (.A(_01244_),
    .X(net2798));
 sky130_fd_sc_hs__buf_2 place2799 (.A(_01236_),
    .X(net2799));
 sky130_fd_sc_hs__buf_1 place2802 (.A(_03004_),
    .X(net2802));
 sky130_fd_sc_hs__buf_1 place2801 (.A(_04110_),
    .X(net2801));
 sky130_fd_sc_hs__buf_1 place2803 (.A(_02989_),
    .X(net2803));
 sky130_fd_sc_hs__buf_1 place2804 (.A(_01218_),
    .X(net2804));
 sky130_fd_sc_hs__bufbuf_8 place2805 (.A(net5090),
    .X(net2805));
 sky130_fd_sc_hs__buf_1 place2806 (.A(_03003_),
    .X(net2806));
 sky130_fd_sc_hs__buf_1 place2807 (.A(_02062_),
    .X(net2807));
 sky130_fd_sc_hs__buf_1 place2809 (.A(_01219_),
    .X(net2809));
 sky130_fd_sc_hs__buf_1 place2811 (.A(net4865),
    .X(net2811));
 sky130_fd_sc_hs__buf_1 place2812 (.A(_05043_),
    .X(net2812));
 sky130_fd_sc_hs__buf_1 place2813 (.A(_05037_),
    .X(net2813));
 sky130_fd_sc_hs__buf_1 place2815 (.A(_05003_),
    .X(net2815));
 sky130_fd_sc_hs__buf_1 place2816 (.A(_04118_),
    .X(net2816));
 sky130_fd_sc_hs__buf_1 place2820 (.A(_05034_),
    .X(net2820));
 sky130_fd_sc_hs__buf_1 place2819 (.A(_05135_),
    .X(net2819));
 sky130_fd_sc_hs__buf_1 place2821 (.A(_05011_),
    .X(net2821));
 sky130_fd_sc_hs__buf_1 place2822 (.A(_05009_),
    .X(net2822));
 sky130_fd_sc_hs__buf_1 place2823 (.A(_05000_),
    .X(net2823));
 sky130_fd_sc_hs__buf_1 place2824 (.A(_04117_),
    .X(net2824));
 sky130_fd_sc_hs__buf_1 place2827 (.A(net2826),
    .X(net2827));
 sky130_fd_sc_hs__buf_1 place2826 (.A(_04111_),
    .X(net2826));
 sky130_fd_sc_hs__buf_1 place2828 (.A(_04108_),
    .X(net2828));
 sky130_fd_sc_hs__buf_1 place2829 (.A(_04106_),
    .X(net2829));
 sky130_fd_sc_hs__buf_1 place2839 (.A(_05027_),
    .X(net2839));
 sky130_fd_sc_hs__buf_1 place2832 (.A(_04104_),
    .X(net2832));
 sky130_fd_sc_hs__buf_1 place2833 (.A(_04078_),
    .X(net2833));
 sky130_fd_sc_hs__buf_1 place2837 (.A(_05094_),
    .X(net2837));
 sky130_fd_sc_hs__buf_1 place2834 (.A(_01249_),
    .X(net2834));
 sky130_fd_sc_hs__buf_2 place2835 (.A(_01105_),
    .X(net2835));
 sky130_fd_sc_hs__buf_1 place2836 (.A(_05134_),
    .X(net2836));
 sky130_fd_sc_hs__buf_2 rebuffer5089 (.A(_05096_),
    .X(net5089));
 sky130_fd_sc_hs__bufbuf_8 place2840 (.A(_04989_),
    .X(net2840));
 sky130_fd_sc_hs__buf_1 place2841 (.A(_04954_),
    .X(net2841));
 sky130_fd_sc_hs__buf_1 place2842 (.A(_04167_),
    .X(net2842));
 sky130_fd_sc_hs__buf_1 place2846 (.A(net2845),
    .X(net2846));
 sky130_fd_sc_hs__buf_1 place2843 (.A(_04137_),
    .X(net2843));
 sky130_fd_sc_hs__buf_1 place2844 (.A(_04116_),
    .X(net2844));
 sky130_fd_sc_hs__buf_2 place2845 (.A(_04101_),
    .X(net2845));
 sky130_fd_sc_hs__buf_1 place2848 (.A(_04077_),
    .X(net2848));
 sky130_fd_sc_hs__buf_1 place2849 (.A(_02987_),
    .X(net2849));
 sky130_fd_sc_hs__bufbuf_8 place2850 (.A(_02984_),
    .X(net2850));
 sky130_fd_sc_hs__buf_1 place2851 (.A(_02970_),
    .X(net2851));
 sky130_fd_sc_hs__buf_1 place2852 (.A(_01235_),
    .X(net2852));
 sky130_fd_sc_hs__buf_1 place2863 (.A(_01397_),
    .X(net2863));
 sky130_fd_sc_hs__buf_1 place2853 (.A(_01210_),
    .X(net2853));
 sky130_fd_sc_hs__bufbuf_8 place2854 (.A(_05047_),
    .X(net2854));
 sky130_fd_sc_hs__bufbuf_8 place2858 (.A(_04194_),
    .X(net2858));
 sky130_fd_sc_hs__buf_4 place2855 (.A(_04988_),
    .X(net2855));
 sky130_fd_sc_hs__buf_1 place2856 (.A(_04953_),
    .X(net2856));
 sky130_fd_sc_hs__bufbuf_8 place2857 (.A(_04236_),
    .X(net2857));
 sky130_fd_sc_hs__buf_1 place2859 (.A(_04166_),
    .X(net2859));
 sky130_fd_sc_hs__buf_1 place2860 (.A(_04136_),
    .X(net2860));
 sky130_fd_sc_hs__buf_1 place2861 (.A(_02959_),
    .X(net2861));
 sky130_fd_sc_hs__buf_1 place2862 (.A(_01397_),
    .X(net2862));
 sky130_fd_sc_hs__buf_1 place2869 (.A(net2868),
    .X(net2869));
 sky130_fd_sc_hs__buf_1 place2864 (.A(_01300_),
    .X(net2864));
 sky130_fd_sc_hs__buf_1 place2865 (.A(_01234_),
    .X(net2865));
 sky130_fd_sc_hs__buf_4 place2868 (.A(_01169_),
    .X(net2868));
 sky130_fd_sc_hs__buf_1 place2866 (.A(_01191_),
    .X(net2866));
 sky130_fd_sc_hs__buf_1 place2867 (.A(_01170_),
    .X(net2867));
 sky130_fd_sc_hs__buf_1 place2870 (.A(_05268_),
    .X(net2870));
 sky130_fd_sc_hs__buf_1 place2873 (.A(_05046_),
    .X(net2873));
 sky130_fd_sc_hs__buf_2 place2874 (.A(_05026_),
    .X(net2874));
 sky130_fd_sc_hs__buf_8 place2877 (.A(_04277_),
    .X(net2877));
 sky130_fd_sc_hs__bufbuf_8 place2876 (.A(_04336_),
    .X(net2876));
 sky130_fd_sc_hs__buf_1 place2881 (.A(_04073_),
    .X(net2881));
 sky130_fd_sc_hs__buf_1 place2885 (.A(_03014_),
    .X(net2885));
 sky130_fd_sc_hs__buf_1 place2886 (.A(_03010_),
    .X(net2886));
 sky130_fd_sc_hs__buf_1 place2887 (.A(_02973_),
    .X(net2887));
 sky130_fd_sc_hs__buf_1 place2889 (.A(_01706_),
    .X(net2889));
 sky130_fd_sc_hs__buf_1 place2892 (.A(_01393_),
    .X(net2892));
 sky130_fd_sc_hs__buf_1 place2893 (.A(_01330_),
    .X(net2893));
 sky130_fd_sc_hs__buf_8 place2894 (.A(_01286_),
    .X(net2894));
 sky130_fd_sc_hs__buf_1 place2897 (.A(net2896),
    .X(net2897));
 sky130_fd_sc_hs__buf_4 place2896 (.A(_01223_),
    .X(net2896));
 sky130_fd_sc_hs__buf_2 place2905 (.A(_04246_),
    .X(net2905));
 sky130_fd_sc_hs__buf_1 place2899 (.A(_01220_),
    .X(net2899));
 sky130_fd_sc_hs__buf_1 place2900 (.A(_01201_),
    .X(net2900));
 sky130_fd_sc_hs__buf_1 place2901 (.A(net4922),
    .X(net2901));
 sky130_fd_sc_hs__buf_1 place2903 (.A(_04951_),
    .X(net2903));
 sky130_fd_sc_hs__buf_1 place2902 (.A(_04984_),
    .X(net2902));
 sky130_fd_sc_hs__buf_1 place2904 (.A(_04307_),
    .X(net2904));
 sky130_fd_sc_hs__buf_2 place2908 (.A(_04081_),
    .X(net2908));
 sky130_fd_sc_hs__buf_4 place2910 (.A(_03118_),
    .X(net2910));
 sky130_fd_sc_hs__buf_1 place2913 (.A(_03013_),
    .X(net2913));
 sky130_fd_sc_hs__buf_1 place2914 (.A(_03001_),
    .X(net2914));
 sky130_fd_sc_hs__buf_1 place2915 (.A(_02983_),
    .X(net2915));
 sky130_fd_sc_hs__bufbuf_8 place2916 (.A(_02974_),
    .X(net2916));
 sky130_fd_sc_hs__buf_1 place2917 (.A(_02362_),
    .X(net2917));
 sky130_fd_sc_hs__buf_4 place2921 (.A(_01429_),
    .X(net2921));
 sky130_fd_sc_hs__buf_1 place2924 (.A(net2923),
    .X(net2924));
 sky130_fd_sc_hs__buf_4 place2923 (.A(_01363_),
    .X(net2923));
 sky130_fd_sc_hs__buf_1 place2927 (.A(net2926),
    .X(net2927));
 sky130_fd_sc_hs__buf_4 place2926 (.A(_01333_),
    .X(net2926));
 sky130_fd_sc_hs__buf_1 place2929 (.A(net2928),
    .X(net2929));
 sky130_fd_sc_hs__buf_4 place2928 (.A(_01303_),
    .X(net2928));
 sky130_fd_sc_hs__buf_1 place2934 (.A(_04982_),
    .X(net2934));
 sky130_fd_sc_hs__buf_1 place2930 (.A(_01200_),
    .X(net2930));
 sky130_fd_sc_hs__buf_1 place2933 (.A(_04996_),
    .X(net2933));
 sky130_fd_sc_hs__bufbuf_8 place2931 (.A(_01152_),
    .X(net2931));
 sky130_fd_sc_hs__buf_2 place2932 (.A(_05005_),
    .X(net2932));
 sky130_fd_sc_hs__bufbuf_8 place2935 (.A(_04950_),
    .X(net2935));
 sky130_fd_sc_hs__buf_1 place2936 (.A(_04133_),
    .X(net2936));
 sky130_fd_sc_hs__buf_1 place2937 (.A(_04068_),
    .X(net2937));
 sky130_fd_sc_hs__buf_1 place2938 (.A(_03148_),
    .X(net2938));
 sky130_fd_sc_hs__buf_1 place2940 (.A(_02939_),
    .X(net2940));
 sky130_fd_sc_hs__buf_1 place2941 (.A(_02481_),
    .X(net2941));
 sky130_fd_sc_hs__buf_1 place2942 (.A(_01151_),
    .X(net2942));
 sky130_fd_sc_hs__buf_2 place2943 (.A(_00993_),
    .X(net2943));
 sky130_fd_sc_hs__buf_1 place2946 (.A(_05509_),
    .X(net2946));
 sky130_fd_sc_hs__buf_2 place2947 (.A(_04995_),
    .X(net2947));
 sky130_fd_sc_hs__buf_1 place2949 (.A(_04949_),
    .X(net2949));
 sky130_fd_sc_hs__buf_1 place2952 (.A(net2951),
    .X(net2952));
 sky130_fd_sc_hs__buf_1 place2950 (.A(_04938_),
    .X(net2950));
 sky130_fd_sc_hs__buf_2 place2951 (.A(_04132_),
    .X(net2951));
 sky130_fd_sc_hs__buf_1 place2953 (.A(_03994_),
    .X(net2953));
 sky130_fd_sc_hs__buf_1 place2954 (.A(_03279_),
    .X(net2954));
 sky130_fd_sc_hs__buf_1 place2959 (.A(_02938_),
    .X(net2959));
 sky130_fd_sc_hs__buf_1 place2960 (.A(_02479_),
    .X(net2960));
 sky130_fd_sc_hs__buf_1 place2961 (.A(net3838),
    .X(net2961));
 sky130_fd_sc_hs__buf_2 place2962 (.A(_01131_),
    .X(net2962));
 sky130_fd_sc_hs__buf_1 place2965 (.A(_00759_),
    .X(net2965));
 sky130_fd_sc_hs__buf_1 place2986 (.A(net2985),
    .X(net2986));
 sky130_fd_sc_hs__buf_1 place2968 (.A(_04994_),
    .X(net2968));
 sky130_fd_sc_hs__buf_1 place2969 (.A(_04990_),
    .X(net2969));
 sky130_fd_sc_hs__buf_1 place2970 (.A(_04987_),
    .X(net2970));
 sky130_fd_sc_hs__buf_1 place2971 (.A(_04983_),
    .X(net2971));
 sky130_fd_sc_hs__buf_1 place2972 (.A(_04978_),
    .X(net2972));
 sky130_fd_sc_hs__buf_1 place2973 (.A(_04965_),
    .X(net2973));
 sky130_fd_sc_hs__buf_1 place2974 (.A(_04948_),
    .X(net2974));
 sky130_fd_sc_hs__buf_2 place2985 (.A(_02927_),
    .X(net2985));
 sky130_fd_sc_hs__buf_1 place2975 (.A(_04895_),
    .X(net2975));
 sky130_fd_sc_hs__buf_2 place2982 (.A(_02980_),
    .X(net2982));
 sky130_fd_sc_hs__bufbuf_8 place2976 (.A(_04131_),
    .X(net2976));
 sky130_fd_sc_hs__buf_1 place2977 (.A(_04074_),
    .X(net2977));
 sky130_fd_sc_hs__buf_1 place2978 (.A(_04043_),
    .X(net2978));
 sky130_fd_sc_hs__bufbuf_8 place2979 (.A(_04026_),
    .X(net2979));
 sky130_fd_sc_hs__buf_1 place2980 (.A(_04021_),
    .X(net2980));
 sky130_fd_sc_hs__buf_1 place2981 (.A(_03443_),
    .X(net2981));
 sky130_fd_sc_hs__buf_2 place2983 (.A(_02964_),
    .X(net2983));
 sky130_fd_sc_hs__buf_4 place2984 (.A(_02956_),
    .X(net2984));
 sky130_fd_sc_hs__buf_1 place2987 (.A(net5123),
    .X(net2987));
 sky130_fd_sc_hs__buf_2 place2988 (.A(_02876_),
    .X(net2988));
 sky130_fd_sc_hs__bufbuf_8 place2990 (.A(_02868_),
    .X(net2990));
 sky130_fd_sc_hs__buf_1 place2991 (.A(_02351_),
    .X(net2991));
 sky130_fd_sc_hs__buf_1 place2993 (.A(_01188_),
    .X(net2993));
 sky130_fd_sc_hs__buf_1 place2994 (.A(_01163_),
    .X(net2994));
 sky130_fd_sc_hs__buf_1 place2995 (.A(net4868),
    .X(net2995));
 sky130_fd_sc_hs__bufbuf_8 place2996 (.A(_01130_),
    .X(net2996));
 sky130_fd_sc_hs__bufbuf_8 place2997 (.A(_01085_),
    .X(net2997));
 sky130_fd_sc_hs__bufbuf_8 place2998 (.A(_01022_),
    .X(net2998));
 sky130_fd_sc_hs__buf_1 place2999 (.A(_00845_),
    .X(net2999));
 sky130_fd_sc_hs__buf_1 place3000 (.A(_05617_),
    .X(net3000));
 sky130_fd_sc_hs__bufbuf_8 place3002 (.A(_05017_),
    .X(net3002));
 sky130_fd_sc_hs__buf_4 place3003 (.A(_05015_),
    .X(net3003));
 sky130_fd_sc_hs__buf_1 place3005 (.A(_04986_),
    .X(net3005));
 sky130_fd_sc_hs__buf_1 place3007 (.A(_04977_),
    .X(net3007));
 sky130_fd_sc_hs__buf_1 place3008 (.A(_04970_),
    .X(net3008));
 sky130_fd_sc_hs__buf_1 place3009 (.A(_04964_),
    .X(net3009));
 sky130_fd_sc_hs__bufbuf_8 place3010 (.A(_04962_),
    .X(net3010));
 sky130_fd_sc_hs__buf_1 place3012 (.A(_04933_),
    .X(net3012));
 sky130_fd_sc_hs__buf_1 place3013 (.A(_04915_),
    .X(net3013));
 sky130_fd_sc_hs__buf_1 place3014 (.A(net5063),
    .X(net3014));
 sky130_fd_sc_hs__buf_1 place3015 (.A(net5096),
    .X(net3015));
 sky130_fd_sc_hs__buf_2 place3016 (.A(_04085_),
    .X(net3016));
 sky130_fd_sc_hs__buf_1 place3018 (.A(_04049_),
    .X(net3018));
 sky130_fd_sc_hs__buf_1 place3019 (.A(net4899),
    .X(net3019));
 sky130_fd_sc_hs__buf_1 place3020 (.A(_04034_),
    .X(net3020));
 sky130_fd_sc_hs__buf_1 place3021 (.A(_04025_),
    .X(net3021));
 sky130_fd_sc_hs__buf_1 place3022 (.A(_04017_),
    .X(net3022));
 sky130_fd_sc_hs__buf_1 place3047 (.A(net3046),
    .X(net3047));
 sky130_fd_sc_hs__clkbuf_2 place3037 (.A(net3036),
    .X(net3037));
 sky130_fd_sc_hs__buf_1 place3026 (.A(_03982_),
    .X(net3026));
 sky130_fd_sc_hs__buf_1 place3029 (.A(_02880_),
    .X(net3029));
 sky130_fd_sc_hs__buf_1 place3027 (.A(_02963_),
    .X(net3027));
 sky130_fd_sc_hs__buf_1 place3028 (.A(_02960_),
    .X(net3028));
 sky130_fd_sc_hs__buf_1 place3030 (.A(_01193_),
    .X(net3030));
 sky130_fd_sc_hs__buf_1 place3031 (.A(_01187_),
    .X(net3031));
 sky130_fd_sc_hs__buf_1 place3032 (.A(_01161_),
    .X(net3032));
 sky130_fd_sc_hs__buf_1 place3033 (.A(_01153_),
    .X(net3033));
 sky130_fd_sc_hs__buf_1 place3034 (.A(_01146_),
    .X(net3034));
 sky130_fd_sc_hs__buf_1 place3035 (.A(_01126_),
    .X(net3035));
 sky130_fd_sc_hs__buf_1 place3036 (.A(_01108_),
    .X(net3036));
 sky130_fd_sc_hs__buf_1 place3038 (.A(_01103_),
    .X(net3038));
 sky130_fd_sc_hs__bufbuf_8 place3039 (.A(_01101_),
    .X(net3039));
 sky130_fd_sc_hs__buf_1 place3040 (.A(_01052_),
    .X(net3040));
 sky130_fd_sc_hs__buf_1 place3041 (.A(_01021_),
    .X(net3041));
 sky130_fd_sc_hs__buf_1 place3042 (.A(_01008_),
    .X(net3042));
 sky130_fd_sc_hs__buf_1 place3043 (.A(_00992_),
    .X(net3043));
 sky130_fd_sc_hs__buf_1 place3044 (.A(_00893_),
    .X(net3044));
 sky130_fd_sc_hs__buf_1 place3045 (.A(net3790),
    .X(net3045));
 sky130_fd_sc_hs__buf_1 place3046 (.A(_00797_),
    .X(net3046));
 sky130_fd_sc_hs__buf_1 place3050 (.A(_04968_),
    .X(net3050));
 sky130_fd_sc_hs__bufbuf_8 place3048 (.A(_05019_),
    .X(net3048));
 sky130_fd_sc_hs__buf_2 place3049 (.A(_05014_),
    .X(net3049));
 sky130_fd_sc_hs__buf_1 place3051 (.A(_04961_),
    .X(net3051));
 sky130_fd_sc_hs__buf_1 place3052 (.A(_04937_),
    .X(net3052));
 sky130_fd_sc_hs__buf_1 place3054 (.A(_04900_),
    .X(net3054));
 sky130_fd_sc_hs__bufbuf_8 place3055 (.A(_04894_),
    .X(net3055));
 sky130_fd_sc_hs__buf_2 place3056 (.A(_04884_),
    .X(net3056));
 sky130_fd_sc_hs__buf_1 place3057 (.A(_04882_),
    .X(net3057));
 sky130_fd_sc_hs__buf_1 place3058 (.A(_04872_),
    .X(net3058));
 sky130_fd_sc_hs__buf_1 place3090 (.A(net3089),
    .X(net3090));
 sky130_fd_sc_hs__buf_1 place3089 (.A(_02232_),
    .X(net3089));
 sky130_fd_sc_hs__buf_1 place3075 (.A(_03924_),
    .X(net3075));
 sky130_fd_sc_hs__buf_1 place3068 (.A(_04020_),
    .X(net3068));
 sky130_fd_sc_hs__buf_4 place3063 (.A(_04084_),
    .X(net3063));
 sky130_fd_sc_hs__bufbuf_8 place3064 (.A(_04070_),
    .X(net3064));
 sky130_fd_sc_hs__bufbuf_8 place3065 (.A(_04069_),
    .X(net3065));
 sky130_fd_sc_hs__bufbuf_8 place3066 (.A(_04024_),
    .X(net3066));
 sky130_fd_sc_hs__buf_1 place3067 (.A(_04020_),
    .X(net3067));
 sky130_fd_sc_hs__buf_1 place3072 (.A(net3071),
    .X(net3072));
 sky130_fd_sc_hs__buf_1 place3069 (.A(_04016_),
    .X(net3069));
 sky130_fd_sc_hs__buf_1 place3070 (.A(_04008_),
    .X(net3070));
 sky130_fd_sc_hs__buf_2 place3071 (.A(_03992_),
    .X(net3071));
 sky130_fd_sc_hs__buf_1 place3074 (.A(net3073),
    .X(net3074));
 sky130_fd_sc_hs__buf_1 place3073 (.A(_03924_),
    .X(net3073));
 sky130_fd_sc_hs__buf_1 place3083 (.A(net3082),
    .X(net3083));
 sky130_fd_sc_hs__buf_1 place3080 (.A(_02924_),
    .X(net3080));
 sky130_fd_sc_hs__bufbuf_8 place3076 (.A(_02953_),
    .X(net3076));
 sky130_fd_sc_hs__bufbuf_8 place3077 (.A(_02948_),
    .X(net3077));
 sky130_fd_sc_hs__buf_1 place3078 (.A(_02942_),
    .X(net3078));
 sky130_fd_sc_hs__bufbuf_8 place3079 (.A(_02937_),
    .X(net3079));
 sky130_fd_sc_hs__buf_1 place3081 (.A(_02886_),
    .X(net3081));
 sky130_fd_sc_hs__buf_2 place3082 (.A(_02883_),
    .X(net3082));
 sky130_fd_sc_hs__buf_1 place3088 (.A(net3086),
    .X(net3088));
 sky130_fd_sc_hs__buf_1 place3084 (.A(_02881_),
    .X(net3084));
 sky130_fd_sc_hs__buf_1 place3087 (.A(net3086),
    .X(net3087));
 sky130_fd_sc_hs__buf_1 place3085 (.A(_02866_),
    .X(net3085));
 sky130_fd_sc_hs__buf_2 place3086 (.A(_02232_),
    .X(net3086));
 sky130_fd_sc_hs__buf_1 place3110 (.A(net3109),
    .X(net3110));
 sky130_fd_sc_hs__buf_1 place3109 (.A(_04871_),
    .X(net3109));
 sky130_fd_sc_hs__buf_1 place3091 (.A(_01192_),
    .X(net3091));
 sky130_fd_sc_hs__buf_1 place3108 (.A(net3106),
    .X(net3108));
 sky130_fd_sc_hs__buf_1 place3102 (.A(net3101),
    .X(net3102));
 sky130_fd_sc_hs__buf_1 place3093 (.A(_00991_),
    .X(net3093));
 sky130_fd_sc_hs__buf_1 place3092 (.A(_01135_),
    .X(net3092));
 sky130_fd_sc_hs__buf_1 place3094 (.A(_00942_),
    .X(net3094));
 sky130_fd_sc_hs__bufbuf_8 place3095 (.A(_04980_),
    .X(net3095));
 sky130_fd_sc_hs__bufbuf_8 place3096 (.A(_04979_),
    .X(net3096));
 sky130_fd_sc_hs__buf_1 place3097 (.A(_04956_),
    .X(net3097));
 sky130_fd_sc_hs__bufbuf_8 place3098 (.A(_04945_),
    .X(net3098));
 sky130_fd_sc_hs__buf_1 place3099 (.A(_04943_),
    .X(net3099));
 sky130_fd_sc_hs__buf_1 place3100 (.A(net5081),
    .X(net3100));
 sky130_fd_sc_hs__buf_1 place3101 (.A(_04936_),
    .X(net3101));
 sky130_fd_sc_hs__buf_1 place3107 (.A(net3106),
    .X(net3107));
 sky130_fd_sc_hs__buf_1 place3103 (.A(_04923_),
    .X(net3103));
 sky130_fd_sc_hs__buf_1 place3104 (.A(_04919_),
    .X(net3104));
 sky130_fd_sc_hs__buf_1 place3105 (.A(_04899_),
    .X(net3105));
 sky130_fd_sc_hs__buf_1 place3106 (.A(_04871_),
    .X(net3106));
 sky130_fd_sc_hs__buf_1 place3116 (.A(net3115),
    .X(net3116));
 sky130_fd_sc_hs__buf_1 place3111 (.A(net5057),
    .X(net3111));
 sky130_fd_sc_hs__bufbuf_8 place3112 (.A(_04083_),
    .X(net3112));
 sky130_fd_sc_hs__buf_1 place3113 (.A(_04056_),
    .X(net3113));
 sky130_fd_sc_hs__buf_1 place3114 (.A(_04045_),
    .X(net3114));
 sky130_fd_sc_hs__buf_2 place3115 (.A(_04030_),
    .X(net3115));
 sky130_fd_sc_hs__buf_1 place3117 (.A(_04023_),
    .X(net3117));
 sky130_fd_sc_hs__buf_1 place3118 (.A(_04019_),
    .X(net3118));
 sky130_fd_sc_hs__buf_1 place3123 (.A(net3122),
    .X(net3123));
 sky130_fd_sc_hs__bufbuf_8 place3119 (.A(_03991_),
    .X(net3119));
 sky130_fd_sc_hs__buf_1 place3120 (.A(_03976_),
    .X(net3120));
 sky130_fd_sc_hs__bufbuf_8 place3121 (.A(_03945_),
    .X(net3121));
 sky130_fd_sc_hs__buf_4 place3122 (.A(_02978_),
    .X(net3122));
 sky130_fd_sc_hs__bufbuf_8 place3124 (.A(_02952_),
    .X(net3124));
 sky130_fd_sc_hs__buf_1 place3125 (.A(_02936_),
    .X(net3125));
 sky130_fd_sc_hs__buf_1 place3126 (.A(_02931_),
    .X(net3126));
 sky130_fd_sc_hs__buf_1 place3130 (.A(_02865_),
    .X(net3130));
 sky130_fd_sc_hs__buf_1 place3127 (.A(_02923_),
    .X(net3127));
 sky130_fd_sc_hs__buf_1 place3128 (.A(_02885_),
    .X(net3128));
 sky130_fd_sc_hs__buf_1 place3129 (.A(_02872_),
    .X(net3129));
 sky130_fd_sc_hs__buf_2 place3131 (.A(_02230_),
    .X(net3131));
 sky130_fd_sc_hs__buf_1 place3140 (.A(net3139),
    .X(net3140));
 sky130_fd_sc_hs__buf_1 place3133 (.A(_01158_),
    .X(net3133));
 sky130_fd_sc_hs__buf_1 place3134 (.A(_01133_),
    .X(net3134));
 sky130_fd_sc_hs__buf_1 place3135 (.A(_01132_),
    .X(net3135));
 sky130_fd_sc_hs__buf_8 place3136 (.A(_01097_),
    .X(net3136));
 sky130_fd_sc_hs__buf_1 place3137 (.A(_01033_),
    .X(net3137));
 sky130_fd_sc_hs__buf_1 place3138 (.A(_00982_),
    .X(net3138));
 sky130_fd_sc_hs__buf_4 place3139 (.A(_00968_),
    .X(net3139));
 sky130_fd_sc_hs__buf_1 place3141 (.A(_00941_),
    .X(net3141));
 sky130_fd_sc_hs__buf_1 place3142 (.A(_00937_),
    .X(net3142));
 sky130_fd_sc_hs__buf_1 place3143 (.A(net4921),
    .X(net3143));
 sky130_fd_sc_hs__buf_1 place3144 (.A(_00902_),
    .X(net3144));
 sky130_fd_sc_hs__buf_1 place3145 (.A(_05013_),
    .X(net3145));
 sky130_fd_sc_hs__bufbuf_8 place3146 (.A(_04971_),
    .X(net3146));
 sky130_fd_sc_hs__buf_1 place3147 (.A(_04934_),
    .X(net3147));
 sky130_fd_sc_hs__buf_1 place3148 (.A(_04925_),
    .X(net3148));
 sky130_fd_sc_hs__bufbuf_8 place3149 (.A(_04921_),
    .X(net3149));
 sky130_fd_sc_hs__buf_1 place3150 (.A(_04917_),
    .X(net3150));
 sky130_fd_sc_hs__buf_1 place3151 (.A(_04909_),
    .X(net3151));
 sky130_fd_sc_hs__buf_1 place3153 (.A(_04883_),
    .X(net3153));
 sky130_fd_sc_hs__buf_1 place3152 (.A(_04892_),
    .X(net3152));
 sky130_fd_sc_hs__buf_4 place3154 (.A(_04880_),
    .X(net3154));
 sky130_fd_sc_hs__bufbuf_8 place3155 (.A(_04086_),
    .X(net3155));
 sky130_fd_sc_hs__bufbuf_8 place3156 (.A(_04082_),
    .X(net3156));
 sky130_fd_sc_hs__buf_1 place3157 (.A(_04058_),
    .X(net3157));
 sky130_fd_sc_hs__buf_1 place3158 (.A(_04053_),
    .X(net3158));
 sky130_fd_sc_hs__bufbuf_8 place3168 (.A(_02965_),
    .X(net3168));
 sky130_fd_sc_hs__buf_1 place3167 (.A(net3166),
    .X(net3167));
 sky130_fd_sc_hs__buf_1 place3160 (.A(_04018_),
    .X(net3160));
 sky130_fd_sc_hs__buf_1 place3161 (.A(net4888),
    .X(net3161));
 sky130_fd_sc_hs__bufbuf_8 place3162 (.A(_04005_),
    .X(net3162));
 sky130_fd_sc_hs__buf_2 place3166 (.A(_02977_),
    .X(net3166));
 sky130_fd_sc_hs__bufbuf_8 place3163 (.A(_03970_),
    .X(net3163));
 sky130_fd_sc_hs__bufbuf_8 place3164 (.A(_03957_),
    .X(net3164));
 sky130_fd_sc_hs__buf_1 place3165 (.A(_03944_),
    .X(net3165));
 sky130_fd_sc_hs__buf_2 place3169 (.A(_02962_),
    .X(net3169));
 sky130_fd_sc_hs__buf_1 place3171 (.A(_02947_),
    .X(net3171));
 sky130_fd_sc_hs__buf_1 place3173 (.A(_02935_),
    .X(net3173));
 sky130_fd_sc_hs__buf_1 place3174 (.A(_02934_),
    .X(net3174));
 sky130_fd_sc_hs__bufbuf_8 place3175 (.A(_02930_),
    .X(net3175));
 sky130_fd_sc_hs__bufbuf_8 place3176 (.A(_02922_),
    .X(net3176));
 sky130_fd_sc_hs__buf_1 place3177 (.A(_02895_),
    .X(net3177));
 sky130_fd_sc_hs__buf_1 place3178 (.A(_02871_),
    .X(net3178));
 sky130_fd_sc_hs__bufbuf_8 place3180 (.A(_01143_),
    .X(net3180));
 sky130_fd_sc_hs__bufbuf_8 place3181 (.A(_01096_),
    .X(net3181));
 sky130_fd_sc_hs__buf_2 place3182 (.A(_01095_),
    .X(net3182));
 sky130_fd_sc_hs__bufbuf_8 place3186 (.A(_00988_),
    .X(net3186));
 sky130_fd_sc_hs__buf_1 place3187 (.A(_00966_),
    .X(net3187));
 sky130_fd_sc_hs__buf_1 place3189 (.A(_00919_),
    .X(net3189));
 sky130_fd_sc_hs__buf_1 place3190 (.A(_00885_),
    .X(net3190));
 sky130_fd_sc_hs__buf_1 place3193 (.A(_00787_),
    .X(net3193));
 sky130_fd_sc_hs__buf_1 place3194 (.A(_04940_),
    .X(net3194));
 sky130_fd_sc_hs__buf_2 place3195 (.A(_04920_),
    .X(net3195));
 sky130_fd_sc_hs__buf_1 place3196 (.A(_04918_),
    .X(net3196));
 sky130_fd_sc_hs__buf_1 place3197 (.A(_04914_),
    .X(net3197));
 sky130_fd_sc_hs__buf_2 place3198 (.A(_04890_),
    .X(net3198));
 sky130_fd_sc_hs__buf_1 place3199 (.A(net5042),
    .X(net3199));
 sky130_fd_sc_hs__buf_1 place3200 (.A(_04869_),
    .X(net3200));
 sky130_fd_sc_hs__bufbuf_8 place3201 (.A(_04057_),
    .X(net3201));
 sky130_fd_sc_hs__bufbuf_8 place3202 (.A(_04052_),
    .X(net3202));
 sky130_fd_sc_hs__buf_1 place3203 (.A(_04047_),
    .X(net3203));
 sky130_fd_sc_hs__buf_1 place3206 (.A(net3205),
    .X(net3206));
 sky130_fd_sc_hs__buf_1 place3204 (.A(_04040_),
    .X(net3204));
 sky130_fd_sc_hs__clkbuf_4 place3205 (.A(_04039_),
    .X(net3205));
 sky130_fd_sc_hs__buf_1 place3207 (.A(_03987_),
    .X(net3207));
 sky130_fd_sc_hs__buf_1 place3224 (.A(_01142_),
    .X(net3224));
 sky130_fd_sc_hs__buf_1 place3215 (.A(_02929_),
    .X(net3215));
 sky130_fd_sc_hs__bufbuf_8 place3208 (.A(_03986_),
    .X(net3208));
 sky130_fd_sc_hs__bufbuf_8 place3209 (.A(_03980_),
    .X(net3209));
 sky130_fd_sc_hs__buf_1 place3210 (.A(_03959_),
    .X(net3210));
 sky130_fd_sc_hs__buf_1 place3211 (.A(_03956_),
    .X(net3211));
 sky130_fd_sc_hs__buf_1 place3212 (.A(_03920_),
    .X(net3212));
 sky130_fd_sc_hs__buf_1 place3214 (.A(_02929_),
    .X(net3214));
 sky130_fd_sc_hs__buf_1 place3213 (.A(_02961_),
    .X(net3213));
 sky130_fd_sc_hs__buf_1 place3216 (.A(_02921_),
    .X(net3216));
 sky130_fd_sc_hs__buf_1 place3217 (.A(_02911_),
    .X(net3217));
 sky130_fd_sc_hs__buf_1 place3219 (.A(net3218),
    .X(net3219));
 sky130_fd_sc_hs__buf_1 place3218 (.A(_02899_),
    .X(net3218));
 sky130_fd_sc_hs__buf_1 place3220 (.A(_02897_),
    .X(net3220));
 sky130_fd_sc_hs__buf_1 place3221 (.A(_02888_),
    .X(net3221));
 sky130_fd_sc_hs__buf_1 place3222 (.A(net5203),
    .X(net3222));
 sky130_fd_sc_hs__bufbuf_8 place3223 (.A(_02863_),
    .X(net3223));
 sky130_fd_sc_hs__bufbuf_8 place3225 (.A(_01137_),
    .X(net3225));
 sky130_fd_sc_hs__buf_2 place3226 (.A(net3801),
    .X(net3226));
 sky130_fd_sc_hs__buf_1 place3227 (.A(_00967_),
    .X(net3227));
 sky130_fd_sc_hs__buf_1 place3229 (.A(net4869),
    .X(net3229));
 sky130_fd_sc_hs__buf_1 place3231 (.A(_00925_),
    .X(net3231));
 sky130_fd_sc_hs__bufbuf_8 place3230 (.A(_00925_),
    .X(net3230));
 sky130_fd_sc_hs__buf_1 place3236 (.A(_00782_),
    .X(net3236));
 sky130_fd_sc_hs__buf_1 place3232 (.A(net4933),
    .X(net3232));
 sky130_fd_sc_hs__buf_1 place3233 (.A(_00898_),
    .X(net3233));
 sky130_fd_sc_hs__bufbuf_8 place3234 (.A(_00877_),
    .X(net3234));
 sky130_fd_sc_hs__buf_1 place3235 (.A(_00860_),
    .X(net3235));
 sky130_fd_sc_hs__buf_4 place3237 (.A(_00733_),
    .X(net3237));
 sky130_fd_sc_hs__buf_1 place3239 (.A(_04922_),
    .X(net3239));
 sky130_fd_sc_hs__buf_2 place3240 (.A(_04913_),
    .X(net3240));
 sky130_fd_sc_hs__buf_1 place3241 (.A(_04911_),
    .X(net3241));
 sky130_fd_sc_hs__buf_1 place3242 (.A(_04906_),
    .X(net3242));
 sky130_fd_sc_hs__buf_1 place3243 (.A(_04878_),
    .X(net3243));
 sky130_fd_sc_hs__buf_4 place3244 (.A(_04867_),
    .X(net3244));
 sky130_fd_sc_hs__buf_2 place3246 (.A(_04833_),
    .X(net3246));
 sky130_fd_sc_hs__buf_1 place3248 (.A(net4891),
    .X(net3248));
 sky130_fd_sc_hs__buf_2 place3249 (.A(_03985_),
    .X(net3249));
 sky130_fd_sc_hs__buf_1 place3252 (.A(net3251),
    .X(net3252));
 sky130_fd_sc_hs__buf_1 place3250 (.A(_03974_),
    .X(net3250));
 sky130_fd_sc_hs__buf_2 place3251 (.A(_03966_),
    .X(net3251));
 sky130_fd_sc_hs__buf_1 place3253 (.A(_03961_),
    .X(net3253));
 sky130_fd_sc_hs__buf_1 place3259 (.A(net3258),
    .X(net3259));
 sky130_fd_sc_hs__buf_1 place3255 (.A(_03958_),
    .X(net3255));
 sky130_fd_sc_hs__buf_1 place3256 (.A(_03913_),
    .X(net3256));
 sky130_fd_sc_hs__bufbuf_8 place3257 (.A(_02954_),
    .X(net3257));
 sky130_fd_sc_hs__buf_2 place3258 (.A(_02925_),
    .X(net3258));
 sky130_fd_sc_hs__buf_1 place3264 (.A(_02869_),
    .X(net3264));
 sky130_fd_sc_hs__bufbuf_8 place3260 (.A(_02919_),
    .X(net3260));
 sky130_fd_sc_hs__buf_1 place3261 (.A(_02917_),
    .X(net3261));
 sky130_fd_sc_hs__bufbuf_8 place3262 (.A(_02908_),
    .X(net3262));
 sky130_fd_sc_hs__buf_1 place3263 (.A(_02892_),
    .X(net3263));
 sky130_fd_sc_hs__bufbuf_8 place3265 (.A(_02862_),
    .X(net3265));
 sky130_fd_sc_hs__buf_1 place3266 (.A(_02199_),
    .X(net3266));
 sky130_fd_sc_hs__buf_1 place3267 (.A(_01028_),
    .X(net3267));
 sky130_fd_sc_hs__buf_1 place3268 (.A(_00984_),
    .X(net3268));
 sky130_fd_sc_hs__buf_1 place3269 (.A(_00961_),
    .X(net3269));
 sky130_fd_sc_hs__bufbuf_8 place3270 (.A(_00917_),
    .X(net3270));
 sky130_fd_sc_hs__buf_1 place3271 (.A(_00817_),
    .X(net3271));
 sky130_fd_sc_hs__buf_1 place3272 (.A(_00781_),
    .X(net3272));
 sky130_fd_sc_hs__buf_1 place3277 (.A(_04912_),
    .X(net3277));
 sky130_fd_sc_hs__bufbuf_8 place3275 (.A(_04974_),
    .X(net3275));
 sky130_fd_sc_hs__buf_1 place3276 (.A(_04912_),
    .X(net3276));
 sky130_fd_sc_hs__buf_1 place3280 (.A(net3279),
    .X(net3280));
 sky130_fd_sc_hs__buf_1 place3279 (.A(net5056),
    .X(net3279));
 sky130_fd_sc_hs__buf_1 place3281 (.A(_04887_),
    .X(net3281));
 sky130_fd_sc_hs__buf_4 place3282 (.A(_04860_),
    .X(net3282));
 sky130_fd_sc_hs__bufbuf_8 place3283 (.A(_04037_),
    .X(net3283));
 sky130_fd_sc_hs__buf_1 place3284 (.A(_03971_),
    .X(net3284));
 sky130_fd_sc_hs__buf_1 place3285 (.A(_03968_),
    .X(net3285));
 sky130_fd_sc_hs__bufbuf_8 place3286 (.A(_03965_),
    .X(net3286));
 sky130_fd_sc_hs__buf_1 place3287 (.A(_03954_),
    .X(net3287));
 sky130_fd_sc_hs__buf_1 place3288 (.A(_03950_),
    .X(net3288));
 sky130_fd_sc_hs__buf_4 place3289 (.A(_03912_),
    .X(net3289));
 sky130_fd_sc_hs__buf_1 place3291 (.A(_03885_),
    .X(net3291));
 sky130_fd_sc_hs__buf_1 place3292 (.A(_03757_),
    .X(net3292));
 sky130_fd_sc_hs__buf_1 place3293 (.A(_02918_),
    .X(net3293));
 sky130_fd_sc_hs__bufbuf_8 place3294 (.A(_02914_),
    .X(net3294));
 sky130_fd_sc_hs__buf_1 place3295 (.A(_02907_),
    .X(net3295));
 sky130_fd_sc_hs__buf_1 place3299 (.A(_02861_),
    .X(net3299));
 sky130_fd_sc_hs__buf_2 place3297 (.A(_02900_),
    .X(net3297));
 sky130_fd_sc_hs__buf_1 place3298 (.A(_02891_),
    .X(net3298));
 sky130_fd_sc_hs__buf_1 place3300 (.A(_02392_),
    .X(net3300));
 sky130_fd_sc_hs__buf_8 place3301 (.A(_02197_),
    .X(net3301));
 sky130_fd_sc_hs__buf_2 place3302 (.A(_01073_),
    .X(net3302));
 sky130_fd_sc_hs__buf_1 place3304 (.A(_00998_),
    .X(net3304));
 sky130_fd_sc_hs__buf_1 place3307 (.A(_00916_),
    .X(net3307));
 sky130_fd_sc_hs__buf_1 place3308 (.A(_00910_),
    .X(net3308));
 sky130_fd_sc_hs__buf_1 place3309 (.A(_00871_),
    .X(net3309));
 sky130_fd_sc_hs__buf_1 place3313 (.A(_00816_),
    .X(net3313));
 sky130_fd_sc_hs__buf_1 place3318 (.A(net3317),
    .X(net3318));
 sky130_fd_sc_hs__buf_1 place3315 (.A(_00779_),
    .X(net3315));
 sky130_fd_sc_hs__buf_1 place3316 (.A(_00611_),
    .X(net3316));
 sky130_fd_sc_hs__buf_2 place3317 (.A(_04908_),
    .X(net3317));
 sky130_fd_sc_hs__buf_1 place3319 (.A(_04903_),
    .X(net3319));
 sky130_fd_sc_hs__buf_1 place3326 (.A(_03963_),
    .X(net3326));
 sky130_fd_sc_hs__buf_1 place3323 (.A(net3321),
    .X(net3323));
 sky130_fd_sc_hs__buf_1 place3322 (.A(net3321),
    .X(net3322));
 sky130_fd_sc_hs__buf_2 place3321 (.A(_04003_),
    .X(net3321));
 sky130_fd_sc_hs__buf_1 place3324 (.A(_03973_),
    .X(net3324));
 sky130_fd_sc_hs__buf_1 place3325 (.A(_03963_),
    .X(net3325));
 sky130_fd_sc_hs__buf_1 place3327 (.A(_03953_),
    .X(net3327));
 sky130_fd_sc_hs__buf_2 place3328 (.A(_03938_),
    .X(net3328));
 sky130_fd_sc_hs__buf_1 place3342 (.A(_00985_),
    .X(net3342));
 sky130_fd_sc_hs__bufbuf_8 place3329 (.A(_03884_),
    .X(net3329));
 sky130_fd_sc_hs__buf_1 place3330 (.A(_03878_),
    .X(net3330));
 sky130_fd_sc_hs__buf_1 place3331 (.A(_03754_),
    .X(net3331));
 sky130_fd_sc_hs__buf_1 place3332 (.A(_02920_),
    .X(net3332));
 sky130_fd_sc_hs__buf_1 place3333 (.A(_02916_),
    .X(net3333));
 sky130_fd_sc_hs__bufbuf_8 place3334 (.A(_02913_),
    .X(net3334));
 sky130_fd_sc_hs__buf_1 place3335 (.A(_02890_),
    .X(net3335));
 sky130_fd_sc_hs__bufbuf_8 place3336 (.A(_02860_),
    .X(net3336));
 sky130_fd_sc_hs__buf_1 place3340 (.A(_01011_),
    .X(net3340));
 sky130_fd_sc_hs__buf_1 place3337 (.A(_02196_),
    .X(net3337));
 sky130_fd_sc_hs__buf_4 place3338 (.A(_02175_),
    .X(net3338));
 sky130_fd_sc_hs__buf_8 place3339 (.A(_01090_),
    .X(net3339));
 sky130_fd_sc_hs__buf_1 place3341 (.A(_00997_),
    .X(net3341));
 sky130_fd_sc_hs__buf_1 place3343 (.A(net4877),
    .X(net3343));
 sky130_fd_sc_hs__buf_1 place3351 (.A(_00837_),
    .X(net3351));
 sky130_fd_sc_hs__bufbuf_8 place3346 (.A(_00926_),
    .X(net3346));
 sky130_fd_sc_hs__buf_1 place3345 (.A(_00962_),
    .X(net3345));
 sky130_fd_sc_hs__buf_1 place3347 (.A(_00920_),
    .X(net3347));
 sky130_fd_sc_hs__bufbuf_8 place3348 (.A(_00874_),
    .X(net3348));
 sky130_fd_sc_hs__buf_1 place3349 (.A(_00856_),
    .X(net3349));
 sky130_fd_sc_hs__buf_1 place3350 (.A(_00837_),
    .X(net3350));
 sky130_fd_sc_hs__buf_1 place3352 (.A(_00832_),
    .X(net3352));
 sky130_fd_sc_hs__buf_2 place3353 (.A(_00786_),
    .X(net3353));
 sky130_fd_sc_hs__buf_2 place3356 (.A(_00737_),
    .X(net3356));
 sky130_fd_sc_hs__bufbuf_8 place3358 (.A(_00732_),
    .X(net3358));
 sky130_fd_sc_hs__buf_1 place3359 (.A(_00724_),
    .X(net3359));
 sky130_fd_sc_hs__buf_1 place3362 (.A(_00152_),
    .X(net3362));
 sky130_fd_sc_hs__buf_1 place3360 (.A(_00710_),
    .X(net3360));
 sky130_fd_sc_hs__buf_1 place3361 (.A(_00680_),
    .X(net3361));
 sky130_fd_sc_hs__bufbuf_8 place3363 (.A(_04973_),
    .X(net3363));
 sky130_fd_sc_hs__buf_1 place3364 (.A(_04958_),
    .X(net3364));
 sky130_fd_sc_hs__buf_1 place3365 (.A(_04904_),
    .X(net3365));
 sky130_fd_sc_hs__buf_1 place3366 (.A(_04875_),
    .X(net3366));
 sky130_fd_sc_hs__buf_1 place3367 (.A(_04865_),
    .X(net3367));
 sky130_fd_sc_hs__buf_1 place3369 (.A(_04863_),
    .X(net3369));
 sky130_fd_sc_hs__buf_1 place3377 (.A(_03883_),
    .X(net3377));
 sky130_fd_sc_hs__bufbuf_8 place3370 (.A(_04849_),
    .X(net3370));
 sky130_fd_sc_hs__buf_1 place3371 (.A(net5061),
    .X(net3371));
 sky130_fd_sc_hs__buf_1 place3375 (.A(_03932_),
    .X(net3375));
 sky130_fd_sc_hs__buf_1 place3372 (.A(_04001_),
    .X(net3372));
 sky130_fd_sc_hs__bufbuf_8 place3373 (.A(_03952_),
    .X(net3373));
 sky130_fd_sc_hs__buf_1 place3374 (.A(_03948_),
    .X(net3374));
 sky130_fd_sc_hs__buf_1 place3376 (.A(_03883_),
    .X(net3376));
 sky130_fd_sc_hs__bufbuf_8 place3378 (.A(_03880_),
    .X(net3378));
 sky130_fd_sc_hs__buf_1 place3379 (.A(_03752_),
    .X(net3379));
 sky130_fd_sc_hs__buf_1 place3381 (.A(_02950_),
    .X(net3381));
 sky130_fd_sc_hs__buf_1 place3382 (.A(_02902_),
    .X(net3382));
 sky130_fd_sc_hs__buf_1 place3383 (.A(_02857_),
    .X(net3383));
 sky130_fd_sc_hs__buf_1 place3387 (.A(_02207_),
    .X(net3387));
 sky130_fd_sc_hs__buf_1 place3386 (.A(_02318_),
    .X(net3386));
 sky130_fd_sc_hs__bufbuf_8 place3390 (.A(_01140_),
    .X(net3390));
 sky130_fd_sc_hs__bufbuf_8 place3395 (.A(_00868_),
    .X(net3395));
 sky130_fd_sc_hs__buf_1 place3391 (.A(_01044_),
    .X(net3391));
 sky130_fd_sc_hs__bufbuf_8 place3392 (.A(_00996_),
    .X(net3392));
 sky130_fd_sc_hs__buf_1 place3393 (.A(_00946_),
    .X(net3393));
 sky130_fd_sc_hs__buf_1 place3394 (.A(_00868_),
    .X(net3394));
 sky130_fd_sc_hs__buf_1 place3396 (.A(_00862_),
    .X(net3396));
 sky130_fd_sc_hs__buf_1 place3397 (.A(_00855_),
    .X(net3397));
 sky130_fd_sc_hs__buf_1 place3399 (.A(_00824_),
    .X(net3399));
 sky130_fd_sc_hs__buf_1 place3403 (.A(_00785_),
    .X(net3403));
 sky130_fd_sc_hs__buf_1 place3405 (.A(_00744_),
    .X(net3405));
 sky130_fd_sc_hs__buf_4 place3406 (.A(_00736_),
    .X(net3406));
 sky130_fd_sc_hs__buf_1 place3410 (.A(net4876),
    .X(net3410));
 sky130_fd_sc_hs__buf_4 place3411 (.A(_00723_),
    .X(net3411));
 sky130_fd_sc_hs__buf_1 place3414 (.A(_00696_),
    .X(net3414));
 sky130_fd_sc_hs__buf_1 place3419 (.A(_00679_),
    .X(net3419));
 sky130_fd_sc_hs__buf_1 place3420 (.A(_00672_),
    .X(net3420));
 sky130_fd_sc_hs__buf_1 place3422 (.A(_04957_),
    .X(net3422));
 sky130_fd_sc_hs__buf_1 place3424 (.A(_04861_),
    .X(net3424));
 sky130_fd_sc_hs__buf_1 place3444 (.A(_02856_),
    .X(net3444));
 sky130_fd_sc_hs__bufbuf_8 place3425 (.A(_04854_),
    .X(net3425));
 sky130_fd_sc_hs__buf_1 place3440 (.A(net3439),
    .X(net3440));
 sky130_fd_sc_hs__bufbuf_8 place3426 (.A(_04848_),
    .X(net3426));
 sky130_fd_sc_hs__bufbuf_8 place3437 (.A(_03908_),
    .X(net3437));
 sky130_fd_sc_hs__bufbuf_8 place3427 (.A(_04835_),
    .X(net3427));
 sky130_fd_sc_hs__buf_1 place3428 (.A(net5086),
    .X(net3428));
 sky130_fd_sc_hs__buf_1 place3430 (.A(_04819_),
    .X(net3430));
 sky130_fd_sc_hs__buf_1 place3429 (.A(_04820_),
    .X(net3429));
 sky130_fd_sc_hs__buf_1 place3431 (.A(_04007_),
    .X(net3431));
 sky130_fd_sc_hs__buf_1 place3432 (.A(_04004_),
    .X(net3432));
 sky130_fd_sc_hs__bufbuf_8 place3433 (.A(_03940_),
    .X(net3433));
 sky130_fd_sc_hs__bufbuf_8 place3434 (.A(_03931_),
    .X(net3434));
 sky130_fd_sc_hs__buf_1 place3435 (.A(_03919_),
    .X(net3435));
 sky130_fd_sc_hs__buf_1 place3436 (.A(_03916_),
    .X(net3436));
 sky130_fd_sc_hs__buf_1 place3438 (.A(_03903_),
    .X(net3438));
 sky130_fd_sc_hs__buf_2 place3439 (.A(_03895_),
    .X(net3439));
 sky130_fd_sc_hs__buf_1 place3441 (.A(_03882_),
    .X(net3441));
 sky130_fd_sc_hs__bufbuf_8 place3442 (.A(_03879_),
    .X(net3442));
 sky130_fd_sc_hs__buf_1 place3443 (.A(_02904_),
    .X(net3443));
 sky130_fd_sc_hs__bufbuf_8 place3445 (.A(_02214_),
    .X(net3445));
 sky130_fd_sc_hs__buf_1 place3446 (.A(_02211_),
    .X(net3446));
 sky130_fd_sc_hs__buf_1 place3452 (.A(_01088_),
    .X(net3452));
 sky130_fd_sc_hs__buf_1 place3447 (.A(_02194_),
    .X(net3447));
 sky130_fd_sc_hs__buf_1 place3450 (.A(_01114_),
    .X(net3450));
 sky130_fd_sc_hs__bufbuf_8 place3448 (.A(_01118_),
    .X(net3448));
 sky130_fd_sc_hs__buf_1 place3449 (.A(_01114_),
    .X(net3449));
 sky130_fd_sc_hs__buf_1 place3451 (.A(_01092_),
    .X(net3451));
 sky130_fd_sc_hs__bufbuf_8 place3457 (.A(_01000_),
    .X(net3457));
 sky130_fd_sc_hs__buf_1 place3463 (.A(_00835_),
    .X(net3463));
 sky130_fd_sc_hs__bufbuf_8 place3460 (.A(_00875_),
    .X(net3460));
 sky130_fd_sc_hs__buf_1 place3461 (.A(_00851_),
    .X(net3461));
 sky130_fd_sc_hs__buf_1 place3462 (.A(_00849_),
    .X(net3462));
 sky130_fd_sc_hs__buf_1 place3464 (.A(_00834_),
    .X(net3464));
 sky130_fd_sc_hs__buf_1 place3471 (.A(_00778_),
    .X(net3471));
 sky130_fd_sc_hs__buf_1 place3466 (.A(_00827_),
    .X(net3466));
 sky130_fd_sc_hs__buf_1 place3467 (.A(_00826_),
    .X(net3467));
 sky130_fd_sc_hs__buf_1 place3468 (.A(_00806_),
    .X(net3468));
 sky130_fd_sc_hs__buf_1 place3469 (.A(_00805_),
    .X(net3469));
 sky130_fd_sc_hs__buf_1 place3470 (.A(_00784_),
    .X(net3470));
 sky130_fd_sc_hs__bufbuf_8 place3472 (.A(_00749_),
    .X(net3472));
 sky130_fd_sc_hs__bufbuf_8 place3473 (.A(_00743_),
    .X(net3473));
 sky130_fd_sc_hs__bufbuf_8 place3474 (.A(_00742_),
    .X(net3474));
 sky130_fd_sc_hs__buf_1 place3475 (.A(_00741_),
    .X(net3475));
 sky130_fd_sc_hs__buf_1 place3476 (.A(_00740_),
    .X(net3476));
 sky130_fd_sc_hs__buf_1 place3477 (.A(_00730_),
    .X(net3477));
 sky130_fd_sc_hs__buf_1 place3479 (.A(_00713_),
    .X(net3479));
 sky130_fd_sc_hs__buf_1 place3481 (.A(_00711_),
    .X(net3481));
 sky130_fd_sc_hs__buf_2 place3487 (.A(_00689_),
    .X(net3487));
 sky130_fd_sc_hs__buf_1 place3488 (.A(_00686_),
    .X(net3488));
 sky130_fd_sc_hs__buf_1 place3492 (.A(net3491),
    .X(net3492));
 sky130_fd_sc_hs__buf_1 place3490 (.A(_00685_),
    .X(net3490));
 sky130_fd_sc_hs__buf_2 place3491 (.A(_00682_),
    .X(net3491));
 sky130_fd_sc_hs__buf_1 place3495 (.A(_00670_),
    .X(net3495));
 sky130_fd_sc_hs__buf_1 place3497 (.A(_00229_),
    .X(net3497));
 sky130_fd_sc_hs__buf_1 place3498 (.A(_00228_),
    .X(net3498));
 sky130_fd_sc_hs__buf_1 place3499 (.A(_00227_),
    .X(net3499));
 sky130_fd_sc_hs__buf_1 place3500 (.A(_00226_),
    .X(net3500));
 sky130_fd_sc_hs__buf_1 place3502 (.A(_00218_),
    .X(net3502));
 sky130_fd_sc_hs__buf_1 place3503 (.A(_00149_),
    .X(net3503));
 sky130_fd_sc_hs__buf_1 place3504 (.A(_00148_),
    .X(net3504));
 sky130_fd_sc_hs__buf_1 place3505 (.A(_00146_),
    .X(net3505));
 sky130_fd_sc_hs__buf_1 place3509 (.A(_00140_),
    .X(net3509));
 sky130_fd_sc_hs__buf_1 place3510 (.A(_00139_),
    .X(net3510));
 sky130_fd_sc_hs__buf_1 place3516 (.A(_00132_),
    .X(net3516));
 sky130_fd_sc_hs__buf_1 place3512 (.A(net3789),
    .X(net3512));
 sky130_fd_sc_hs__buf_1 place3515 (.A(net3514),
    .X(net3515));
 sky130_fd_sc_hs__buf_1 place3513 (.A(_00134_),
    .X(net3513));
 sky130_fd_sc_hs__buf_4 place3514 (.A(_00133_),
    .X(net3514));
 sky130_fd_sc_hs__buf_1 place3517 (.A(_00131_),
    .X(net3517));
 sky130_fd_sc_hs__buf_1 place3518 (.A(_00130_),
    .X(net3518));
 sky130_fd_sc_hs__buf_1 place3519 (.A(_00129_),
    .X(net3519));
 sky130_fd_sc_hs__buf_1 place3523 (.A(_00127_),
    .X(net3523));
 sky130_fd_sc_hs__buf_8 place3528 (.A(_00124_),
    .X(net3528));
 sky130_fd_sc_hs__buf_4 place3530 (.A(_00122_),
    .X(net3530));
 sky130_fd_sc_hs__buf_1 place3532 (.A(_00121_),
    .X(net3532));
 sky130_fd_sc_hs__clkbuf_2 place3535 (.A(_00118_),
    .X(net3535));
 sky130_fd_sc_hs__buf_1 place3537 (.A(_00117_),
    .X(net3537));
 sky130_fd_sc_hs__buf_1 place3540 (.A(_00114_),
    .X(net3540));
 sky130_fd_sc_hs__buf_2 place3541 (.A(_00112_),
    .X(net3541));
 sky130_fd_sc_hs__buf_1 place3543 (.A(_00111_),
    .X(net3543));
 sky130_fd_sc_hs__buf_1 place3545 (.A(_00109_),
    .X(net3545));
 sky130_fd_sc_hs__buf_1 place3547 (.A(_00107_),
    .X(net3547));
 sky130_fd_sc_hs__buf_1 place3550 (.A(_00105_),
    .X(net3550));
 sky130_fd_sc_hs__buf_1 place3552 (.A(_00103_),
    .X(net3552));
 sky130_fd_sc_hs__buf_1 place3554 (.A(_00101_),
    .X(net3554));
 sky130_fd_sc_hs__buf_1 place3556 (.A(_00099_),
    .X(net3556));
 sky130_fd_sc_hs__buf_1 place3558 (.A(_00097_),
    .X(net3558));
 sky130_fd_sc_hs__buf_1 place3560 (.A(_00095_),
    .X(net3560));
 sky130_fd_sc_hs__buf_1 place3562 (.A(_00092_),
    .X(net3562));
 sky130_fd_sc_hs__buf_1 place3572 (.A(_04817_),
    .X(net3572));
 sky130_fd_sc_hs__buf_1 place3564 (.A(_00090_),
    .X(net3564));
 sky130_fd_sc_hs__bufbuf_8 place3565 (.A(_04843_),
    .X(net3565));
 sky130_fd_sc_hs__buf_1 place3566 (.A(_04839_),
    .X(net3566));
 sky130_fd_sc_hs__buf_1 place3570 (.A(net3569),
    .X(net3570));
 sky130_fd_sc_hs__buf_1 place3567 (.A(_04830_),
    .X(net3567));
 sky130_fd_sc_hs__buf_1 place3568 (.A(_04825_),
    .X(net3568));
 sky130_fd_sc_hs__buf_1 place3569 (.A(_04824_),
    .X(net3569));
 sky130_fd_sc_hs__buf_1 place3571 (.A(_04817_),
    .X(net3571));
 sky130_fd_sc_hs__bufbuf_8 place3574 (.A(_03989_),
    .X(net3574));
 sky130_fd_sc_hs__buf_1 place3573 (.A(_04009_),
    .X(net3573));
 sky130_fd_sc_hs__buf_1 place3575 (.A(_03984_),
    .X(net3575));
 sky130_fd_sc_hs__buf_1 place3576 (.A(_03951_),
    .X(net3576));
 sky130_fd_sc_hs__bufbuf_8 place3578 (.A(_03935_),
    .X(net3578));
 sky130_fd_sc_hs__bufbuf_8 place3579 (.A(_03934_),
    .X(net3579));
 sky130_fd_sc_hs__bufbuf_8 place3581 (.A(_03930_),
    .X(net3581));
 sky130_fd_sc_hs__buf_1 place3582 (.A(_03929_),
    .X(net3582));
 sky130_fd_sc_hs__buf_1 place3583 (.A(_03918_),
    .X(net3583));
 sky130_fd_sc_hs__buf_1 place3584 (.A(_03917_),
    .X(net3584));
 sky130_fd_sc_hs__buf_1 place3585 (.A(_03915_),
    .X(net3585));
 sky130_fd_sc_hs__buf_1 place3609 (.A(_00210_),
    .X(net3609));
 sky130_fd_sc_hs__buf_1 place3587 (.A(_03914_),
    .X(net3587));
 sky130_fd_sc_hs__buf_1 place3588 (.A(_03909_),
    .X(net3588));
 sky130_fd_sc_hs__bufbuf_8 place3589 (.A(_03907_),
    .X(net3589));
 sky130_fd_sc_hs__bufbuf_8 place3590 (.A(_03901_),
    .X(net3590));
 sky130_fd_sc_hs__bufbuf_8 place3591 (.A(_03898_),
    .X(net3591));
 sky130_fd_sc_hs__bufbuf_8 place3592 (.A(_03897_),
    .X(net3592));
 sky130_fd_sc_hs__buf_1 place3593 (.A(_03894_),
    .X(net3593));
 sky130_fd_sc_hs__bufbuf_8 place3594 (.A(_03893_),
    .X(net3594));
 sky130_fd_sc_hs__bufbuf_8 place3595 (.A(_03892_),
    .X(net3595));
 sky130_fd_sc_hs__buf_1 place3596 (.A(_03891_),
    .X(net3596));
 sky130_fd_sc_hs__bufbuf_8 place3597 (.A(_03889_),
    .X(net3597));
 sky130_fd_sc_hs__buf_1 place3598 (.A(_03888_),
    .X(net3598));
 sky130_fd_sc_hs__bufbuf_8 place3605 (.A(_03872_),
    .X(net3605));
 sky130_fd_sc_hs__buf_1 place3600 (.A(_03887_),
    .X(net3600));
 sky130_fd_sc_hs__buf_1 place3599 (.A(_03887_),
    .X(net3599));
 sky130_fd_sc_hs__bufbuf_8 place3601 (.A(_03886_),
    .X(net3601));
 sky130_fd_sc_hs__buf_1 place3602 (.A(_03875_),
    .X(net3602));
 sky130_fd_sc_hs__buf_1 place3603 (.A(_03874_),
    .X(net3603));
 sky130_fd_sc_hs__buf_1 place3604 (.A(_03872_),
    .X(net3604));
 sky130_fd_sc_hs__bufbuf_8 place3606 (.A(_02903_),
    .X(net3606));
 sky130_fd_sc_hs__bufbuf_8 place3607 (.A(_02889_),
    .X(net3607));
 sky130_fd_sc_hs__bufbuf_8 place3608 (.A(_00210_),
    .X(net3608));
 sky130_fd_sc_hs__buf_1 place3610 (.A(_02224_),
    .X(net3610));
 sky130_fd_sc_hs__bufbuf_8 place3611 (.A(_02223_),
    .X(net3611));
 sky130_fd_sc_hs__buf_1 place3612 (.A(_02220_),
    .X(net3612));
 sky130_fd_sc_hs__buf_1 place3614 (.A(_02219_),
    .X(net3614));
 sky130_fd_sc_hs__buf_1 place3615 (.A(_02218_),
    .X(net3615));
 sky130_fd_sc_hs__bufbuf_8 place3616 (.A(_02213_),
    .X(net3616));
 sky130_fd_sc_hs__bufbuf_8 place3617 (.A(_02212_),
    .X(net3617));
 sky130_fd_sc_hs__buf_1 place3618 (.A(_02210_),
    .X(net3618));
 sky130_fd_sc_hs__buf_1 place3619 (.A(_02209_),
    .X(net3619));
 sky130_fd_sc_hs__bufbuf_8 place3620 (.A(_02205_),
    .X(net3620));
 sky130_fd_sc_hs__buf_1 place3622 (.A(_02201_),
    .X(net3622));
 sky130_fd_sc_hs__buf_1 place3624 (.A(_02200_),
    .X(net3624));
 sky130_fd_sc_hs__buf_1 place3625 (.A(_02198_),
    .X(net3625));
 sky130_fd_sc_hs__buf_1 place3626 (.A(_02193_),
    .X(net3626));
 sky130_fd_sc_hs__buf_1 place3628 (.A(_02191_),
    .X(net3628));
 sky130_fd_sc_hs__buf_1 place3629 (.A(_02190_),
    .X(net3629));
 sky130_fd_sc_hs__buf_1 place3630 (.A(_02188_),
    .X(net3630));
 sky130_fd_sc_hs__buf_1 place3633 (.A(_02111_),
    .X(net3633));
 sky130_fd_sc_hs__buf_1 place3631 (.A(_00211_),
    .X(net3631));
 sky130_fd_sc_hs__buf_1 place3632 (.A(_02111_),
    .X(net3632));
 sky130_fd_sc_hs__buf_1 place3635 (.A(_02108_),
    .X(net3635));
 sky130_fd_sc_hs__buf_1 place3634 (.A(_02108_),
    .X(net3634));
 sky130_fd_sc_hs__buf_1 place3640 (.A(_02087_),
    .X(net3640));
 sky130_fd_sc_hs__bufbuf_8 place3637 (.A(_02104_),
    .X(net3637));
 sky130_fd_sc_hs__bufbuf_8 place3638 (.A(_02095_),
    .X(net3638));
 sky130_fd_sc_hs__buf_1 place3639 (.A(_02087_),
    .X(net3639));
 sky130_fd_sc_hs__buf_1 place3642 (.A(_02084_),
    .X(net3642));
 sky130_fd_sc_hs__buf_1 place3641 (.A(_02084_),
    .X(net3641));
 sky130_fd_sc_hs__bufbuf_8 place3644 (.A(_02077_),
    .X(net3644));
 sky130_fd_sc_hs__buf_1 place3643 (.A(_02077_),
    .X(net3643));
 sky130_fd_sc_hs__buf_1 place3647 (.A(_02067_),
    .X(net3647));
 sky130_fd_sc_hs__bufbuf_8 place3645 (.A(_02073_),
    .X(net3645));
 sky130_fd_sc_hs__buf_1 place3646 (.A(_02067_),
    .X(net3646));
 sky130_fd_sc_hs__bufbuf_8 place3648 (.A(_02058_),
    .X(net3648));
 sky130_fd_sc_hs__bufbuf_8 place3649 (.A(_02048_),
    .X(net3649));
 sky130_fd_sc_hs__buf_1 place3654 (.A(_02034_),
    .X(net3654));
 sky130_fd_sc_hs__buf_1 place3652 (.A(_02038_),
    .X(net3652));
 sky130_fd_sc_hs__buf_1 place3651 (.A(_02038_),
    .X(net3651));
 sky130_fd_sc_hs__buf_1 place3653 (.A(_02034_),
    .X(net3653));
 sky130_fd_sc_hs__buf_2 place3657 (.A(_02025_),
    .X(net3657));
 sky130_fd_sc_hs__bufbuf_8 place3655 (.A(_02028_),
    .X(net3655));
 sky130_fd_sc_hs__buf_1 place3656 (.A(_02025_),
    .X(net3656));
 sky130_fd_sc_hs__buf_1 place3660 (.A(net3659),
    .X(net3660));
 sky130_fd_sc_hs__buf_1 place3659 (.A(_02019_),
    .X(net3659));
 sky130_fd_sc_hs__buf_1 place3668 (.A(_01965_),
    .X(net3668));
 sky130_fd_sc_hs__buf_1 place3661 (.A(_02015_),
    .X(net3661));
 sky130_fd_sc_hs__bufbuf_8 place3665 (.A(_01980_),
    .X(net3665));
 sky130_fd_sc_hs__bufbuf_8 place3662 (.A(_02006_),
    .X(net3662));
 sky130_fd_sc_hs__bufbuf_8 place3663 (.A(_01989_),
    .X(net3663));
 sky130_fd_sc_hs__buf_1 place3664 (.A(_01985_),
    .X(net3664));
 sky130_fd_sc_hs__buf_1 place3666 (.A(_01976_),
    .X(net3666));
 sky130_fd_sc_hs__bufbuf_8 place3667 (.A(_01965_),
    .X(net3667));
 sky130_fd_sc_hs__buf_1 place3670 (.A(_01950_),
    .X(net3670));
 sky130_fd_sc_hs__buf_1 place3669 (.A(_01950_),
    .X(net3669));
 sky130_fd_sc_hs__bufbuf_8 place3672 (.A(_00150_),
    .X(net3672));
 sky130_fd_sc_hs__buf_1 place3671 (.A(_00150_),
    .X(net3671));
 sky130_fd_sc_hs__buf_4 place3673 (.A(_00658_),
    .X(net3673));
 sky130_fd_sc_hs__buf_1 place3674 (.A(_00613_),
    .X(net3674));
 sky130_fd_sc_hs__buf_1 place3678 (.A(\u_window_buffer.write_ptr[8] ),
    .X(net3678));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hs__buf_1 place3680 (.A(\u_window_buffer.write_ptr[7] ),
    .X(net3680));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hs__buf_1 place3688 (.A(\u_window_buffer.write_ptr[2] ),
    .X(net3688));
 sky130_fd_sc_hs__buf_1 place3681 (.A(\u_window_buffer.write_ptr[6] ),
    .X(net3681));
 sky130_fd_sc_hs__buf_1 place3682 (.A(\u_window_buffer.write_ptr[5] ),
    .X(net3682));
 sky130_fd_sc_hs__buf_1 place3683 (.A(\u_window_buffer.write_ptr[4] ),
    .X(net3683));
 sky130_fd_sc_hs__buf_1 place3686 (.A(\u_window_buffer.write_ptr[30] ),
    .X(net3686));
 sky130_fd_sc_hs__buf_1 place3685 (.A(\u_window_buffer.write_ptr[31] ),
    .X(net3685));
 sky130_fd_sc_hs__buf_1 place3684 (.A(\u_window_buffer.write_ptr[31] ),
    .X(net3684));
 sky130_fd_sc_hs__buf_1 place3687 (.A(\u_window_buffer.write_ptr[2] ),
    .X(net3687));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hs__buf_1 place3689 (.A(\u_window_buffer.write_ptr[29] ),
    .X(net3689));
 sky130_fd_sc_hs__buf_1 place3690 (.A(\u_window_buffer.write_ptr[28] ),
    .X(net3690));
 sky130_fd_sc_hs__buf_1 place3691 (.A(\u_window_buffer.write_ptr[27] ),
    .X(net3691));
 sky130_fd_sc_hs__buf_1 place3692 (.A(\u_window_buffer.write_ptr[26] ),
    .X(net3692));
 sky130_fd_sc_hs__buf_1 place3693 (.A(\u_window_buffer.write_ptr[25] ),
    .X(net3693));
 sky130_fd_sc_hs__buf_1 place3694 (.A(\u_window_buffer.write_ptr[24] ),
    .X(net3694));
 sky130_fd_sc_hs__buf_1 place3696 (.A(\u_window_buffer.write_ptr[23] ),
    .X(net3696));
 sky130_fd_sc_hs__buf_1 place3695 (.A(\u_window_buffer.write_ptr[23] ),
    .X(net3695));
 sky130_fd_sc_hs__buf_1 place3698 (.A(\u_window_buffer.write_ptr[22] ),
    .X(net3698));
 sky130_fd_sc_hs__buf_1 place3697 (.A(\u_window_buffer.write_ptr[22] ),
    .X(net3697));
 sky130_fd_sc_hs__buf_1 place3700 (.A(\u_window_buffer.write_ptr[21] ),
    .X(net3700));
 sky130_fd_sc_hs__buf_1 place3699 (.A(\u_window_buffer.write_ptr[21] ),
    .X(net3699));
 sky130_fd_sc_hs__buf_4 place3783 (.A(net3782),
    .X(net3783));
 sky130_fd_sc_hs__buf_1 place3701 (.A(\u_window_buffer.write_ptr[20] ),
    .X(net3701));
 sky130_fd_sc_hs__buf_1 place3702 (.A(\u_window_buffer.write_ptr[1] ),
    .X(net3702));
 sky130_fd_sc_hs__buf_1 place3725 (.A(\u_window_buffer.read_ptr[28] ),
    .X(net3725));
 sky130_fd_sc_hs__buf_1 place3703 (.A(\u_window_buffer.write_ptr[19] ),
    .X(net3703));
 sky130_fd_sc_hs__buf_1 place3704 (.A(\u_window_buffer.write_ptr[18] ),
    .X(net3704));
 sky130_fd_sc_hs__buf_1 place3705 (.A(\u_window_buffer.write_ptr[17] ),
    .X(net3705));
 sky130_fd_sc_hs__buf_1 place3706 (.A(\u_window_buffer.write_ptr[16] ),
    .X(net3706));
 sky130_fd_sc_hs__buf_1 place3707 (.A(\u_window_buffer.write_ptr[15] ),
    .X(net3707));
 sky130_fd_sc_hs__buf_1 place3708 (.A(\u_window_buffer.write_ptr[14] ),
    .X(net3708));
 sky130_fd_sc_hs__buf_1 place3709 (.A(\u_window_buffer.write_ptr[13] ),
    .X(net3709));
 sky130_fd_sc_hs__buf_1 place3710 (.A(\u_window_buffer.write_ptr[12] ),
    .X(net3710));
 sky130_fd_sc_hs__buf_1 place3711 (.A(\u_window_buffer.write_ptr[11] ),
    .X(net3711));
 sky130_fd_sc_hs__buf_1 place3712 (.A(\u_window_buffer.write_ptr[10] ),
    .X(net3712));
 sky130_fd_sc_hs__buf_1 place3713 (.A(net5075),
    .X(net3713));
 sky130_fd_sc_hs__buf_1 place3714 (.A(\u_window_buffer.read_ptr[9] ),
    .X(net3714));
 sky130_fd_sc_hs__buf_1 place3715 (.A(\u_window_buffer.read_ptr[8] ),
    .X(net3715));
 sky130_fd_sc_hs__buf_1 place3716 (.A(\u_window_buffer.read_ptr[7] ),
    .X(net3716));
 sky130_fd_sc_hs__clkbuf_2 place3717 (.A(\u_window_buffer.read_ptr[6] ),
    .X(net3717));
 sky130_fd_sc_hs__clkbuf_4 place3718 (.A(\u_window_buffer.read_ptr[5] ),
    .X(net3718));
 sky130_fd_sc_hs__buf_2 place3719 (.A(\u_window_buffer.read_ptr[4] ),
    .X(net3719));
 sky130_fd_sc_hs__clkbuf_2 place3720 (.A(\u_window_buffer.read_ptr[3] ),
    .X(net3720));
 sky130_fd_sc_hs__buf_1 place3721 (.A(\u_window_buffer.read_ptr[31] ),
    .X(net3721));
 sky130_fd_sc_hs__buf_1 place3722 (.A(\u_window_buffer.read_ptr[30] ),
    .X(net3722));
 sky130_fd_sc_hs__clkbuf_2 place3723 (.A(\u_window_buffer.read_ptr[2] ),
    .X(net3723));
 sky130_fd_sc_hs__buf_1 place3724 (.A(\u_window_buffer.read_ptr[29] ),
    .X(net3724));
 sky130_fd_sc_hs__buf_1 place3726 (.A(\u_window_buffer.read_ptr[27] ),
    .X(net3726));
 sky130_fd_sc_hs__buf_1 place3727 (.A(\u_window_buffer.read_ptr[26] ),
    .X(net3727));
 sky130_fd_sc_hs__buf_1 place3728 (.A(\u_window_buffer.read_ptr[25] ),
    .X(net3728));
 sky130_fd_sc_hs__buf_1 place3729 (.A(\u_window_buffer.read_ptr[24] ),
    .X(net3729));
 sky130_fd_sc_hs__buf_1 place3730 (.A(\u_window_buffer.read_ptr[23] ),
    .X(net3730));
 sky130_fd_sc_hs__buf_1 place3731 (.A(\u_window_buffer.read_ptr[22] ),
    .X(net3731));
 sky130_fd_sc_hs__buf_1 place3732 (.A(\u_window_buffer.read_ptr[21] ),
    .X(net3732));
 sky130_fd_sc_hs__buf_1 place3733 (.A(\u_window_buffer.read_ptr[20] ),
    .X(net3733));
 sky130_fd_sc_hs__buf_4 place3782 (.A(_05774_),
    .X(net3782));
 sky130_fd_sc_hs__buf_1 place3734 (.A(\u_window_buffer.read_ptr[19] ),
    .X(net3734));
 sky130_fd_sc_hs__buf_1 place3735 (.A(\u_window_buffer.read_ptr[18] ),
    .X(net3735));
 sky130_fd_sc_hs__buf_1 place3736 (.A(\u_window_buffer.read_ptr[17] ),
    .X(net3736));
 sky130_fd_sc_hs__buf_1 place3737 (.A(\u_window_buffer.read_ptr[16] ),
    .X(net3737));
 sky130_fd_sc_hs__buf_1 place3738 (.A(\u_window_buffer.read_ptr[15] ),
    .X(net3738));
 sky130_fd_sc_hs__buf_1 place3739 (.A(\u_window_buffer.read_ptr[14] ),
    .X(net3739));
 sky130_fd_sc_hs__clkbuf_2 place3740 (.A(\u_window_buffer.read_ptr[13] ),
    .X(net3740));
 sky130_fd_sc_hs__buf_1 place3741 (.A(\u_window_buffer.read_ptr[12] ),
    .X(net3741));
 sky130_fd_sc_hs__buf_1 place3742 (.A(\u_window_buffer.read_ptr[11] ),
    .X(net3742));
 sky130_fd_sc_hs__clkbuf_2 place3743 (.A(\u_window_buffer.read_ptr[10] ),
    .X(net3743));
 sky130_fd_sc_hs__buf_2 place3744 (.A(\u_window_buffer.read_ptr[0] ),
    .X(net3744));
 sky130_fd_sc_hs__buf_4 place3781 (.A(_05774_),
    .X(net3781));
 sky130_fd_sc_hs__clkbuf_2 place3745 (.A(\u_window_buffer.internal_read_ptr[9] ),
    .X(net3745));
 sky130_fd_sc_hs__buf_1 place3773 (.A(net3772),
    .X(net3773));
 sky130_fd_sc_hs__clkbuf_4 place3746 (.A(\u_window_buffer.internal_read_ptr[8] ),
    .X(net3746));
 sky130_fd_sc_hs__buf_4 place3747 (.A(\u_window_buffer.internal_read_ptr[7] ),
    .X(net3747));
 sky130_fd_sc_hs__clkbuf_8 place3748 (.A(\u_window_buffer.internal_read_ptr[6] ),
    .X(net3748));
 sky130_fd_sc_hs__buf_8 place3749 (.A(\u_window_buffer.internal_read_ptr[5] ),
    .X(net3749));
 sky130_fd_sc_hs__clkbuf_2 place3750 (.A(\u_window_buffer.internal_read_ptr[4] ),
    .X(net3750));
 sky130_fd_sc_hs__buf_1 place3751 (.A(\u_window_buffer.internal_read_ptr[3] ),
    .X(net3751));
 sky130_fd_sc_hs__buf_1 place3752 (.A(\u_window_buffer.internal_read_ptr[31] ),
    .X(net3752));
 sky130_fd_sc_hs__buf_1 place3753 (.A(\u_window_buffer.internal_read_ptr[30] ),
    .X(net3753));
 sky130_fd_sc_hs__buf_1 place3754 (.A(\u_window_buffer.internal_read_ptr[2] ),
    .X(net3754));
 sky130_fd_sc_hs__buf_1 place3755 (.A(\u_window_buffer.internal_read_ptr[29] ),
    .X(net3755));
 sky130_fd_sc_hs__buf_1 place3756 (.A(\u_window_buffer.internal_read_ptr[28] ),
    .X(net3756));
 sky130_fd_sc_hs__buf_1 place3757 (.A(\u_window_buffer.internal_read_ptr[27] ),
    .X(net3757));
 sky130_fd_sc_hs__buf_1 place3758 (.A(\u_window_buffer.internal_read_ptr[26] ),
    .X(net3758));
 sky130_fd_sc_hs__buf_1 place3759 (.A(\u_window_buffer.internal_read_ptr[25] ),
    .X(net3759));
 sky130_fd_sc_hs__buf_1 place3760 (.A(\u_window_buffer.internal_read_ptr[24] ),
    .X(net3760));
 sky130_fd_sc_hs__buf_1 place3761 (.A(\u_window_buffer.internal_read_ptr[23] ),
    .X(net3761));
 sky130_fd_sc_hs__buf_1 place3762 (.A(\u_window_buffer.internal_read_ptr[22] ),
    .X(net3762));
 sky130_fd_sc_hs__buf_1 place3763 (.A(\u_window_buffer.internal_read_ptr[21] ),
    .X(net3763));
 sky130_fd_sc_hs__buf_1 place3764 (.A(\u_window_buffer.internal_read_ptr[20] ),
    .X(net3764));
 sky130_fd_sc_hs__buf_2 place3765 (.A(\u_window_buffer.internal_read_ptr[1] ),
    .X(net3765));
 sky130_fd_sc_hs__buf_1 place3766 (.A(\u_window_buffer.internal_read_ptr[19] ),
    .X(net3766));
 sky130_fd_sc_hs__clkbuf_2 place3767 (.A(\u_window_buffer.internal_read_ptr[18] ),
    .X(net3767));
 sky130_fd_sc_hs__buf_1 place3768 (.A(\u_window_buffer.internal_read_ptr[17] ),
    .X(net3768));
 sky130_fd_sc_hs__buf_1 place3769 (.A(\u_window_buffer.internal_read_ptr[16] ),
    .X(net3769));
 sky130_fd_sc_hs__buf_1 place3770 (.A(\u_window_buffer.internal_read_ptr[15] ),
    .X(net3770));
 sky130_fd_sc_hs__buf_1 place3771 (.A(\u_window_buffer.internal_read_ptr[14] ),
    .X(net3771));
 sky130_fd_sc_hs__buf_8 place3772 (.A(\u_window_buffer.internal_read_ptr[13] ),
    .X(net3772));
 sky130_fd_sc_hs__buf_1 place3774 (.A(\u_window_buffer.internal_read_ptr[12] ),
    .X(net3774));
 sky130_fd_sc_hs__clkbuf_2 place3775 (.A(\u_window_buffer.internal_read_ptr[11] ),
    .X(net3775));
 sky130_fd_sc_hs__clkbuf_2 place3776 (.A(\u_window_buffer.internal_read_ptr[10] ),
    .X(net3776));
 sky130_fd_sc_hs__buf_2 place3777 (.A(\u_window_buffer.current_state[3] ),
    .X(net3777));
 sky130_fd_sc_hs__buf_4 place3778 (.A(\u_window_buffer.current_state[2] ),
    .X(net3778));
 sky130_fd_sc_hs__buf_1 place3779 (.A(\u_hamming_window.hamming_state[2] ),
    .X(net3779));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hs__buf_4 place3784 (.A(net211),
    .X(net3784));
 sky130_fd_sc_hs__buf_1 place3785 (.A(net3784),
    .X(net3785));
 sky130_fd_sc_hs__buf_16 place1847 (.A(net1845),
    .X(net1847));
 sky130_fd_sc_hs__buf_16 place1853 (.A(net5106),
    .X(net1853));
 sky130_fd_sc_hs__buf_1 place1862 (.A(_05698_),
    .X(net1862));
 sky130_fd_sc_hs__buf_1 place1863 (.A(_05698_),
    .X(net1863));
 sky130_fd_sc_hs__buf_2 place1866 (.A(net3786),
    .X(net1866));
 sky130_fd_sc_hs__buf_1 place1867 (.A(_01963_),
    .X(net1867));
 sky130_fd_sc_hs__buf_1 place1869 (.A(net1868),
    .X(net1869));
 sky130_fd_sc_hs__buf_1 rebuffer5203 (.A(_02870_),
    .X(net5203));
 sky130_fd_sc_hs__buf_16 place1873 (.A(_03688_),
    .X(net1873));
 sky130_fd_sc_hs__buf_1 place1910 (.A(_03670_),
    .X(net1910));
 sky130_fd_sc_hs__buf_1 place1912 (.A(_03657_),
    .X(net1912));
 sky130_fd_sc_hs__buf_1 place1918 (.A(_03669_),
    .X(net1918));
 sky130_fd_sc_hs__buf_1 place1920 (.A(_03658_),
    .X(net1920));
 sky130_fd_sc_hs__buf_1 place1921 (.A(net1920),
    .X(net1921));
 sky130_fd_sc_hs__buf_1 place1926 (.A(_03628_),
    .X(net1926));
 sky130_fd_sc_hs__buf_1 place1927 (.A(_01912_),
    .X(net1927));
 sky130_fd_sc_hs__buf_1 place1946 (.A(net1945),
    .X(net1946));
 sky130_fd_sc_hs__buf_1 place1955 (.A(_04718_),
    .X(net1955));
 sky130_fd_sc_hs__buf_1 place1959 (.A(_03615_),
    .X(net1959));
 sky130_fd_sc_hs__buf_1 place1961 (.A(_05605_),
    .X(net1961));
 sky130_fd_sc_hs__buf_1 place1966 (.A(_04701_),
    .X(net1966));
 sky130_fd_sc_hs__buf_1 place1968 (.A(_01899_),
    .X(net1968));
 sky130_fd_sc_hs__buf_1 place1970 (.A(net1969),
    .X(net1970));
 sky130_fd_sc_hs__buf_1 place1971 (.A(_01845_),
    .X(net1971));
 sky130_fd_sc_hs__buf_1 place1972 (.A(_01845_),
    .X(net1972));
 sky130_fd_sc_hs__buf_1 place1974 (.A(_05618_),
    .X(net1974));
 sky130_fd_sc_hs__buf_1 place1979 (.A(_03644_),
    .X(net1979));
 sky130_fd_sc_hs__buf_1 place1985 (.A(_04704_),
    .X(net1985));
 sky130_fd_sc_hs__buf_1 place1986 (.A(_04690_),
    .X(net1986));
 sky130_fd_sc_hs__buf_1 place1987 (.A(_03606_),
    .X(net1987));
 sky130_fd_sc_hs__buf_1 place1989 (.A(net1988),
    .X(net1989));
 sky130_fd_sc_hs__buf_1 place1996 (.A(_04688_),
    .X(net1996));
 sky130_fd_sc_hs__buf_1 place1997 (.A(net1996),
    .X(net1997));
 sky130_fd_sc_hs__buf_2 place2016 (.A(_05621_),
    .X(net2016));
 sky130_fd_sc_hs__buf_1 place2017 (.A(net2016),
    .X(net2017));
 sky130_fd_sc_hs__buf_2 place2031 (.A(_05549_),
    .X(net2031));
 sky130_fd_sc_hs__buf_1 place2032 (.A(net5083),
    .X(net2032));
 sky130_fd_sc_hs__buf_1 place2033 (.A(_05549_),
    .X(net2033));
 sky130_fd_sc_hs__buf_1 place2039 (.A(net2038),
    .X(net2039));
 sky130_fd_sc_hs__bufbuf_8 place2050 (.A(_04664_),
    .X(net2050));
 sky130_fd_sc_hs__buf_1 place2051 (.A(_01810_),
    .X(net2051));
 sky130_fd_sc_hs__bufbuf_8 place2052 (.A(_04666_),
    .X(net2052));
 sky130_fd_sc_hs__buf_1 place2064 (.A(_04646_),
    .X(net2064));
 sky130_fd_sc_hs__buf_1 place2070 (.A(net5043),
    .X(net2070));
 sky130_fd_sc_hs__buf_2 place2074 (.A(_01771_),
    .X(net2074));
 sky130_fd_sc_hs__buf_1 place2076 (.A(net2075),
    .X(net2076));
 sky130_fd_sc_hs__buf_1 place2077 (.A(net2075),
    .X(net2077));
 sky130_fd_sc_hs__buf_1 place2080 (.A(net4890),
    .X(net2080));
 sky130_fd_sc_hs__buf_1 place2083 (.A(net2082),
    .X(net2083));
 sky130_fd_sc_hs__buf_1 place2085 (.A(net5128),
    .X(net2085));
 sky130_fd_sc_hs__buf_1 place2086 (.A(_01792_),
    .X(net2086));
 sky130_fd_sc_hs__buf_1 place2107 (.A(_05506_),
    .X(net2107));
 sky130_fd_sc_hs__buf_1 place2108 (.A(net2107),
    .X(net2108));
 sky130_fd_sc_hs__buf_1 place2113 (.A(_01745_),
    .X(net2113));
 sky130_fd_sc_hs__buf_1 place2118 (.A(_04602_),
    .X(net2118));
 sky130_fd_sc_hs__buf_1 place2123 (.A(_01778_),
    .X(net2123));
 sky130_fd_sc_hs__buf_1 place2124 (.A(_05511_),
    .X(net2124));
 sky130_fd_sc_hs__buf_1 place2127 (.A(_04588_),
    .X(net2127));
 sky130_fd_sc_hs__buf_2 place2135 (.A(net2134),
    .X(net2135));
 sky130_fd_sc_hs__buf_4 place2136 (.A(net2135),
    .X(net2136));
 sky130_fd_sc_hs__buf_1 place2138 (.A(_03495_),
    .X(net2138));
 sky130_fd_sc_hs__buf_1 place2139 (.A(_03491_),
    .X(net2139));
 sky130_fd_sc_hs__buf_1 place2150 (.A(net2149),
    .X(net2150));
 sky130_fd_sc_hs__buf_1 place2153 (.A(net4906),
    .X(net2153));
 sky130_fd_sc_hs__buf_1 place2174 (.A(_04564_),
    .X(net2174));
 sky130_fd_sc_hs__buf_1 place2175 (.A(_04562_),
    .X(net2175));
 sky130_fd_sc_hs__buf_1 place2188 (.A(_03447_),
    .X(net2188));
 sky130_fd_sc_hs__buf_1 place2192 (.A(net5049),
    .X(net2192));
 sky130_fd_sc_hs__buf_1 place2193 (.A(_04535_),
    .X(net2193));
 sky130_fd_sc_hs__bufbuf_8 place2207 (.A(_01673_),
    .X(net2207));
 sky130_fd_sc_hs__buf_1 place2214 (.A(_03426_),
    .X(net2214));
 sky130_fd_sc_hs__buf_1 place2223 (.A(_04512_),
    .X(net2223));
 sky130_fd_sc_hs__buf_1 place2230 (.A(net2229),
    .X(net2230));
 sky130_fd_sc_hs__buf_1 place2237 (.A(_03395_),
    .X(net2237));
 sky130_fd_sc_hs__buf_1 place2239 (.A(_04516_),
    .X(net2239));
 sky130_fd_sc_hs__buf_1 place2241 (.A(_04493_),
    .X(net2241));
 sky130_fd_sc_hs__buf_1 place2244 (.A(_03420_),
    .X(net2244));
 sky130_fd_sc_hs__buf_1 place2273 (.A(_04471_),
    .X(net2273));
 sky130_fd_sc_hs__buf_1 place2275 (.A(_05381_),
    .X(net2275));
 sky130_fd_sc_hs__bufbuf_8 place2276 (.A(_04468_),
    .X(net2276));
 sky130_fd_sc_hs__buf_1 place2288 (.A(net2287),
    .X(net2288));
 sky130_fd_sc_hs__buf_1 place2305 (.A(_03339_),
    .X(net2305));
 sky130_fd_sc_hs__buf_1 place2313 (.A(_01590_),
    .X(net2313));
 sky130_fd_sc_hs__buf_1 place2314 (.A(_04455_),
    .X(net2314));
 sky130_fd_sc_hs__buf_1 place2316 (.A(_04436_),
    .X(net2316));
 sky130_fd_sc_hs__buf_1 place2321 (.A(_03319_),
    .X(net2321));
 sky130_fd_sc_hs__buf_1 place2349 (.A(_04412_),
    .X(net2349));
 sky130_fd_sc_hs__buf_1 place2350 (.A(_04412_),
    .X(net2350));
 sky130_fd_sc_hs__bufbuf_8 place2355 (.A(_03328_),
    .X(net2355));
 sky130_fd_sc_hs__buf_1 place2357 (.A(_03302_),
    .X(net2357));
 sky130_fd_sc_hs__buf_1 place2359 (.A(_04443_),
    .X(net2359));
 sky130_fd_sc_hs__bufbuf_8 place2367 (.A(_01573_),
    .X(net2367));
 sky130_fd_sc_hs__buf_1 place2372 (.A(_05316_),
    .X(net2372));
 sky130_fd_sc_hs__buf_1 place2373 (.A(_05285_),
    .X(net2373));
 sky130_fd_sc_hs__buf_1 place2374 (.A(_04414_),
    .X(net2374));
 sky130_fd_sc_hs__buf_1 place2377 (.A(net2376),
    .X(net2377));
 sky130_fd_sc_hs__buf_1 place2392 (.A(_04381_),
    .X(net2392));
 sky130_fd_sc_hs__buf_1 place2394 (.A(_03282_),
    .X(net2394));
 sky130_fd_sc_hs__buf_1 place2428 (.A(net5102),
    .X(net2428));
 sky130_fd_sc_hs__buf_1 place2431 (.A(_01490_),
    .X(net2431));
 sky130_fd_sc_hs__buf_1 place2446 (.A(_03231_),
    .X(net2446));
 sky130_fd_sc_hs__buf_1 place2449 (.A(_05247_),
    .X(net2449));
 sky130_fd_sc_hs__buf_1 place2452 (.A(_04350_),
    .X(net2452));
 sky130_fd_sc_hs__buf_1 place2502 (.A(_05230_),
    .X(net2502));
 sky130_fd_sc_hs__buf_1 place2504 (.A(_05210_),
    .X(net2504));
 sky130_fd_sc_hs__buf_1 place2505 (.A(_04303_),
    .X(net2505));
 sky130_fd_sc_hs__buf_1 place2506 (.A(_03208_),
    .X(net2506));
 sky130_fd_sc_hs__buf_2 place2508 (.A(net2507),
    .X(net2508));
 sky130_fd_sc_hs__buf_1 place2514 (.A(_05209_),
    .X(net2514));
 sky130_fd_sc_hs__buf_1 place2517 (.A(_04302_),
    .X(net2517));
 sky130_fd_sc_hs__bufbuf_8 place2537 (.A(_04308_),
    .X(net2537));
 sky130_fd_sc_hs__buf_1 place2545 (.A(_01417_),
    .X(net2545));
 sky130_fd_sc_hs__buf_1 place2582 (.A(_04278_),
    .X(net2582));
 sky130_fd_sc_hs__bufbuf_8 place2591 (.A(_04266_),
    .X(net2591));
 sky130_fd_sc_hs__buf_1 place2639 (.A(_05115_),
    .X(net2639));
 sky130_fd_sc_hs__buf_1 place2650 (.A(_01343_),
    .X(net2650));
 sky130_fd_sc_hs__buf_1 place2654 (.A(_05127_),
    .X(net2654));
 sky130_fd_sc_hs__buf_1 place2655 (.A(_05127_),
    .X(net2655));
 sky130_fd_sc_hs__buf_1 place2665 (.A(_03099_),
    .X(net2665));
 sky130_fd_sc_hs__buf_1 place2668 (.A(_03083_),
    .X(net2668));
 sky130_fd_sc_hs__buf_1 place2677 (.A(net2676),
    .X(net2677));
 sky130_fd_sc_hs__buf_1 place2680 (.A(_01322_),
    .X(net2680));
 sky130_fd_sc_hs__buf_1 place2684 (.A(_05095_),
    .X(net2684));
 sky130_fd_sc_hs__buf_1 place2685 (.A(_05088_),
    .X(net2685));
 sky130_fd_sc_hs__buf_2 place2690 (.A(_01327_),
    .X(net2690));
 sky130_fd_sc_hs__clkbuf_2 place2693 (.A(_05090_),
    .X(net2693));
 sky130_fd_sc_hs__buf_1 place2694 (.A(_05078_),
    .X(net2694));
 sky130_fd_sc_hs__buf_1 place2722 (.A(net2721),
    .X(net2722));
 sky130_fd_sc_hs__buf_1 place2730 (.A(_05070_),
    .X(net2730));
 sky130_fd_sc_hs__bufbuf_8 place2734 (.A(_05069_),
    .X(net2734));
 sky130_fd_sc_hs__buf_1 place2737 (.A(_04156_),
    .X(net2737));
 sky130_fd_sc_hs__buf_1 place2749 (.A(_01261_),
    .X(net2749));
 sky130_fd_sc_hs__buf_1 place2754 (.A(net5193),
    .X(net2754));
 sky130_fd_sc_hs__buf_1 place2759 (.A(net2758),
    .X(net2759));
 sky130_fd_sc_hs__buf_1 place2761 (.A(_03009_),
    .X(net2761));
 sky130_fd_sc_hs__buf_1 place2762 (.A(_01265_),
    .X(net2762));
 sky130_fd_sc_hs__buf_1 place2764 (.A(net2763),
    .X(net2764));
 sky130_fd_sc_hs__buf_1 place2769 (.A(_04125_),
    .X(net2769));
 sky130_fd_sc_hs__buf_1 place2771 (.A(_03008_),
    .X(net2771));
 sky130_fd_sc_hs__buf_1 place2775 (.A(_05059_),
    .X(net2775));
 sky130_fd_sc_hs__buf_2 place2776 (.A(_05038_),
    .X(net2776));
 sky130_fd_sc_hs__buf_1 place2777 (.A(net5070),
    .X(net2777));
 sky130_fd_sc_hs__buf_1 place2778 (.A(_03006_),
    .X(net2778));
 sky130_fd_sc_hs__buf_1 place2779 (.A(net5121),
    .X(net2779));
 sky130_fd_sc_hs__buf_1 place2780 (.A(net4895),
    .X(net2780));
 sky130_fd_sc_hs__buf_1 place2781 (.A(_01230_),
    .X(net2781));
 sky130_fd_sc_hs__buf_1 place2783 (.A(net2782),
    .X(net2783));
 sky130_fd_sc_hs__buf_1 place2786 (.A(net2785),
    .X(net2786));
 sky130_fd_sc_hs__buf_1 place2788 (.A(net2787),
    .X(net2788));
 sky130_fd_sc_hs__buf_1 place2792 (.A(_02996_),
    .X(net2792));
 sky130_fd_sc_hs__buf_1 place2800 (.A(net2799),
    .X(net2800));
 sky130_fd_sc_hs__buf_1 place2808 (.A(_01229_),
    .X(net2808));
 sky130_fd_sc_hs__buf_1 place2810 (.A(_01219_),
    .X(net2810));
 sky130_fd_sc_hs__bufbuf_8 place2814 (.A(_05036_),
    .X(net2814));
 sky130_fd_sc_hs__buf_1 place2817 (.A(_04118_),
    .X(net2817));
 sky130_fd_sc_hs__buf_1 place2818 (.A(_04094_),
    .X(net2818));
 sky130_fd_sc_hs__buf_1 place2825 (.A(_04117_),
    .X(net2825));
 sky130_fd_sc_hs__buf_1 place2830 (.A(net2829),
    .X(net2830));
 sky130_fd_sc_hs__buf_1 place2831 (.A(net2829),
    .X(net2831));
 sky130_fd_sc_hs__buf_1 place2847 (.A(net2845),
    .X(net2847));
 sky130_fd_sc_hs__buf_4 place2871 (.A(_05121_),
    .X(net2871));
 sky130_fd_sc_hs__buf_1 place2872 (.A(net2871),
    .X(net2872));
 sky130_fd_sc_hs__bufbuf_8 place2875 (.A(_04998_),
    .X(net2875));
 sky130_fd_sc_hs__buf_1 place2878 (.A(_04274_),
    .X(net2878));
 sky130_fd_sc_hs__buf_1 place2879 (.A(_04235_),
    .X(net2879));
 sky130_fd_sc_hs__buf_1 place2880 (.A(_04193_),
    .X(net2880));
 sky130_fd_sc_hs__buf_1 place2882 (.A(_03135_),
    .X(net2882));
 sky130_fd_sc_hs__buf_1 place2883 (.A(_03098_),
    .X(net2883));
 sky130_fd_sc_hs__buf_1 place2884 (.A(_03046_),
    .X(net2884));
 sky130_fd_sc_hs__buf_1 place2888 (.A(net5124),
    .X(net2888));
 sky130_fd_sc_hs__buf_1 place2890 (.A(_01679_),
    .X(net2890));
 sky130_fd_sc_hs__buf_1 place2891 (.A(_01396_),
    .X(net2891));
 sky130_fd_sc_hs__buf_1 place2895 (.A(net2894),
    .X(net2895));
 sky130_fd_sc_hs__buf_1 place2898 (.A(net2897),
    .X(net2898));
 sky130_fd_sc_hs__buf_1 place2906 (.A(net2905),
    .X(net2906));
 sky130_fd_sc_hs__bufbuf_8 place2907 (.A(_04134_),
    .X(net2907));
 sky130_fd_sc_hs__buf_1 place2909 (.A(_04072_),
    .X(net2909));
 sky130_fd_sc_hs__buf_1 place2911 (.A(_03072_),
    .X(net2911));
 sky130_fd_sc_hs__buf_1 place2912 (.A(_03045_),
    .X(net2912));
 sky130_fd_sc_hs__buf_1 place2918 (.A(_01638_),
    .X(net2918));
 sky130_fd_sc_hs__buf_1 place2919 (.A(_01494_),
    .X(net2919));
 sky130_fd_sc_hs__buf_4 place2920 (.A(_01460_),
    .X(net2920));
 sky130_fd_sc_hs__buf_1 place2922 (.A(net2921),
    .X(net2922));
 sky130_fd_sc_hs__buf_1 place2925 (.A(net2923),
    .X(net2925));
 sky130_fd_sc_hs__bufbuf_8 place2939 (.A(_02967_),
    .X(net2939));
 sky130_fd_sc_hs__buf_1 place2944 (.A(_00762_),
    .X(net2944));
 sky130_fd_sc_hs__buf_1 place2945 (.A(net2944),
    .X(net2945));
 sky130_fd_sc_hs__buf_1 place2948 (.A(_04981_),
    .X(net2948));
 sky130_fd_sc_hs__bufbuf_8 place2955 (.A(_03070_),
    .X(net2955));
 sky130_fd_sc_hs__bufbuf_8 place2956 (.A(net5170),
    .X(net2956));
 sky130_fd_sc_hs__buf_1 place2957 (.A(_02966_),
    .X(net2957));
 sky130_fd_sc_hs__buf_1 place2958 (.A(net5144),
    .X(net2958));
 sky130_fd_sc_hs__buf_1 place2963 (.A(_01023_),
    .X(net2963));
 sky130_fd_sc_hs__buf_1 place2964 (.A(net4874),
    .X(net2964));
 sky130_fd_sc_hs__buf_4 place2966 (.A(net2965),
    .X(net2966));
 sky130_fd_sc_hs__buf_1 place2967 (.A(_00759_),
    .X(net2967));
 sky130_fd_sc_hs__buf_1 place2989 (.A(net2988),
    .X(net2989));
 sky130_fd_sc_hs__buf_2 place2992 (.A(_01207_),
    .X(net2992));
 sky130_fd_sc_hs__bufbuf_8 place3001 (.A(_05018_),
    .X(net3001));
 sky130_fd_sc_hs__buf_1 place3004 (.A(_04993_),
    .X(net3004));
 sky130_fd_sc_hs__buf_1 place3006 (.A(_04986_),
    .X(net3006));
 sky130_fd_sc_hs__bufbuf_8 place3011 (.A(_04942_),
    .X(net3011));
 sky130_fd_sc_hs__bufbuf_8 place3017 (.A(_04079_),
    .X(net3017));
 sky130_fd_sc_hs__buf_1 place3023 (.A(_03995_),
    .X(net3023));
 sky130_fd_sc_hs__buf_1 place3024 (.A(net3023),
    .X(net3024));
 sky130_fd_sc_hs__buf_1 place3025 (.A(_03995_),
    .X(net3025));
 sky130_fd_sc_hs__bufbuf_8 place3053 (.A(_04932_),
    .X(net3053));
 sky130_fd_sc_hs__buf_1 place3059 (.A(_04872_),
    .X(net3059));
 sky130_fd_sc_hs__buf_1 place3060 (.A(_04872_),
    .X(net3060));
 sky130_fd_sc_hs__buf_1 place3061 (.A(_04872_),
    .X(net3061));
 sky130_fd_sc_hs__buf_1 place3062 (.A(net3061),
    .X(net3062));
 sky130_fd_sc_hs__buf_4 place3132 (.A(net3131),
    .X(net3132));
 sky130_fd_sc_hs__buf_1 place3159 (.A(_04053_),
    .X(net3159));
 sky130_fd_sc_hs__buf_1 place3170 (.A(net3169),
    .X(net3170));
 sky130_fd_sc_hs__buf_1 place3172 (.A(_02947_),
    .X(net3172));
 sky130_fd_sc_hs__buf_1 place3179 (.A(_02864_),
    .X(net3179));
 sky130_fd_sc_hs__buf_1 place3183 (.A(net3182),
    .X(net3183));
 sky130_fd_sc_hs__buf_1 place3184 (.A(_01041_),
    .X(net3184));
 sky130_fd_sc_hs__buf_1 place3185 (.A(_00989_),
    .X(net3185));
 sky130_fd_sc_hs__buf_1 place3188 (.A(_00953_),
    .X(net3188));
 sky130_fd_sc_hs__buf_1 place3191 (.A(_00878_),
    .X(net3191));
 sky130_fd_sc_hs__buf_1 place3192 (.A(_00865_),
    .X(net3192));
 sky130_fd_sc_hs__buf_1 place3228 (.A(_00954_),
    .X(net3228));
 sky130_fd_sc_hs__buf_1 rebuffer5065 (.A(_05039_),
    .X(net5065));
 sky130_fd_sc_hs__buf_1 place3245 (.A(net3244),
    .X(net3245));
 sky130_fd_sc_hs__bufbuf_8 place3247 (.A(_04054_),
    .X(net3247));
 sky130_fd_sc_hs__buf_1 place3254 (.A(net3253),
    .X(net3254));
 sky130_fd_sc_hs__buf_1 place3273 (.A(_00775_),
    .X(net3273));
 sky130_fd_sc_hs__bufbuf_8 place3274 (.A(_00716_),
    .X(net3274));
 sky130_fd_sc_hs__buf_1 place3278 (.A(net3277),
    .X(net3278));
 sky130_fd_sc_hs__buf_1 place3290 (.A(net3289),
    .X(net3290));
 sky130_fd_sc_hs__buf_1 place3296 (.A(_02907_),
    .X(net3296));
 sky130_fd_sc_hs__buf_1 place3303 (.A(net3302),
    .X(net3303));
 sky130_fd_sc_hs__buf_1 place3305 (.A(_00927_),
    .X(net3305));
 sky130_fd_sc_hs__buf_8 place3306 (.A(_00921_),
    .X(net3306));
 sky130_fd_sc_hs__buf_2 place3310 (.A(_00864_),
    .X(net3310));
 sky130_fd_sc_hs__buf_1 place3311 (.A(_00838_),
    .X(net3311));
 sky130_fd_sc_hs__buf_1 place3312 (.A(_00833_),
    .X(net3312));
 sky130_fd_sc_hs__buf_1 place3314 (.A(_00816_),
    .X(net3314));
 sky130_fd_sc_hs__buf_1 place3320 (.A(_04903_),
    .X(net3320));
 sky130_fd_sc_hs__clkbuf_2 place3344 (.A(_00977_),
    .X(net3344));
 sky130_fd_sc_hs__buf_1 place3354 (.A(_00777_),
    .X(net3354));
 sky130_fd_sc_hs__buf_1 place3355 (.A(_00745_),
    .X(net3355));
 sky130_fd_sc_hs__buf_1 place3357 (.A(_00737_),
    .X(net3357));
 sky130_fd_sc_hs__buf_1 place3368 (.A(net3367),
    .X(net3368));
 sky130_fd_sc_hs__buf_1 place3380 (.A(_02976_),
    .X(net3380));
 sky130_fd_sc_hs__buf_1 place3384 (.A(_02852_),
    .X(net3384));
 sky130_fd_sc_hs__buf_1 place3385 (.A(_02852_),
    .X(net3385));
 sky130_fd_sc_hs__bufbuf_8 place3388 (.A(_02203_),
    .X(net3388));
 sky130_fd_sc_hs__buf_1 place3389 (.A(_02195_),
    .X(net3389));
 sky130_fd_sc_hs__buf_1 place3398 (.A(net3791),
    .X(net3398));
 sky130_fd_sc_hs__buf_1 place3400 (.A(_00814_),
    .X(net3400));
 sky130_fd_sc_hs__buf_1 place3401 (.A(_00810_),
    .X(net3401));
 sky130_fd_sc_hs__bufbuf_8 place3402 (.A(_00809_),
    .X(net3402));
 sky130_fd_sc_hs__buf_1 place3404 (.A(_00750_),
    .X(net3404));
 sky130_fd_sc_hs__buf_1 place3407 (.A(net3406),
    .X(net3407));
 sky130_fd_sc_hs__buf_2 place3408 (.A(_00731_),
    .X(net3408));
 sky130_fd_sc_hs__buf_1 place3409 (.A(net3408),
    .X(net3409));
 sky130_fd_sc_hs__buf_1 place3412 (.A(_00719_),
    .X(net3412));
 sky130_fd_sc_hs__buf_1 place3413 (.A(_00715_),
    .X(net3413));
 sky130_fd_sc_hs__bufbuf_8 place3415 (.A(_00691_),
    .X(net3415));
 sky130_fd_sc_hs__buf_1 place3416 (.A(_00687_),
    .X(net3416));
 sky130_fd_sc_hs__buf_1 place3417 (.A(_00683_),
    .X(net3417));
 sky130_fd_sc_hs__buf_1 place3418 (.A(_00683_),
    .X(net3418));
 sky130_fd_sc_hs__buf_1 place3421 (.A(_00214_),
    .X(net3421));
 sky130_fd_sc_hs__buf_1 place3423 (.A(_04862_),
    .X(net3423));
 sky130_fd_sc_hs__bufbuf_8 place3453 (.A(_01075_),
    .X(net3453));
 sky130_fd_sc_hs__buf_1 place3454 (.A(_01070_),
    .X(net3454));
 sky130_fd_sc_hs__bufbuf_8 place3455 (.A(_01043_),
    .X(net3455));
 sky130_fd_sc_hs__buf_1 place3456 (.A(_01037_),
    .X(net3456));
 sky130_fd_sc_hs__buf_1 place3458 (.A(_00995_),
    .X(net3458));
 sky130_fd_sc_hs__buf_1 place3459 (.A(_00911_),
    .X(net3459));
 sky130_fd_sc_hs__buf_1 place3465 (.A(_00834_),
    .X(net3465));
 sky130_fd_sc_hs__buf_1 place3478 (.A(_00714_),
    .X(net3478));
 sky130_fd_sc_hs__buf_4 place3480 (.A(net3479),
    .X(net3480));
 sky130_fd_sc_hs__buf_2 place3482 (.A(_00699_),
    .X(net3482));
 sky130_fd_sc_hs__buf_1 place3483 (.A(_00698_),
    .X(net3483));
 sky130_fd_sc_hs__buf_2 place3484 (.A(_00695_),
    .X(net3484));
 sky130_fd_sc_hs__buf_1 place3485 (.A(net3484),
    .X(net3485));
 sky130_fd_sc_hs__buf_2 place3486 (.A(_00694_),
    .X(net3486));
 sky130_fd_sc_hs__buf_1 place3489 (.A(net3488),
    .X(net3489));
 sky130_fd_sc_hs__buf_2 place3493 (.A(_00681_),
    .X(net3493));
 sky130_fd_sc_hs__buf_1 place3494 (.A(net3493),
    .X(net3494));
 sky130_fd_sc_hs__buf_1 place3496 (.A(net3495),
    .X(net3496));
 sky130_fd_sc_hs__buf_1 place3501 (.A(_00219_),
    .X(net3501));
 sky130_fd_sc_hs__buf_1 place3506 (.A(_00145_),
    .X(net3506));
 sky130_fd_sc_hs__buf_1 place3507 (.A(_00144_),
    .X(net3507));
 sky130_fd_sc_hs__buf_1 place3508 (.A(_00142_),
    .X(net3508));
 sky130_fd_sc_hs__buf_1 place3511 (.A(_00138_),
    .X(net3511));
 sky130_fd_sc_hs__buf_1 place3520 (.A(_00129_),
    .X(net3520));
 sky130_fd_sc_hs__buf_8 place3521 (.A(_00128_),
    .X(net3521));
 sky130_fd_sc_hs__buf_1 place3522 (.A(net3521),
    .X(net3522));
 sky130_fd_sc_hs__buf_1 place3524 (.A(net3523),
    .X(net3524));
 sky130_fd_sc_hs__buf_1 place3525 (.A(_00126_),
    .X(net3525));
 sky130_fd_sc_hs__buf_1 place3526 (.A(_00126_),
    .X(net3526));
 sky130_fd_sc_hs__buf_1 place3527 (.A(_00126_),
    .X(net3527));
 sky130_fd_sc_hs__buf_1 place3529 (.A(net3528),
    .X(net3529));
 sky130_fd_sc_hs__buf_1 place3531 (.A(net3530),
    .X(net3531));
 sky130_fd_sc_hs__clkbuf_2 place3533 (.A(_00120_),
    .X(net3533));
 sky130_fd_sc_hs__buf_1 place3534 (.A(net3533),
    .X(net3534));
 sky130_fd_sc_hs__buf_1 place3536 (.A(net3535),
    .X(net3536));
 sky130_fd_sc_hs__buf_8 place3538 (.A(_00116_),
    .X(net3538));
 sky130_fd_sc_hs__buf_1 place3539 (.A(net3538),
    .X(net3539));
 sky130_fd_sc_hs__buf_1 place3542 (.A(net3541),
    .X(net3542));
 sky130_fd_sc_hs__buf_1 place3544 (.A(_00110_),
    .X(net3544));
 sky130_fd_sc_hs__dlymetal6s2s_1 place3546 (.A(_00108_),
    .X(net3546));
 sky130_fd_sc_hs__buf_2 place3548 (.A(_00106_),
    .X(net3548));
 sky130_fd_sc_hs__buf_1 place3549 (.A(net3548),
    .X(net3549));
 sky130_fd_sc_hs__buf_2 place3551 (.A(_00104_),
    .X(net3551));
 sky130_fd_sc_hs__buf_2 place3553 (.A(_00102_),
    .X(net3553));
 sky130_fd_sc_hs__buf_1 place3555 (.A(_00100_),
    .X(net3555));
 sky130_fd_sc_hs__buf_1 place3557 (.A(_00098_),
    .X(net3557));
 sky130_fd_sc_hs__buf_1 place3559 (.A(_00096_),
    .X(net3559));
 sky130_fd_sc_hs__buf_1 place3561 (.A(_00094_),
    .X(net3561));
 sky130_fd_sc_hs__buf_1 place3563 (.A(_00092_),
    .X(net3563));
 sky130_fd_sc_hs__bufbuf_8 place3577 (.A(_03939_),
    .X(net3577));
 sky130_fd_sc_hs__buf_1 place3580 (.A(_03933_),
    .X(net3580));
 sky130_fd_sc_hs__buf_1 place3586 (.A(_03915_),
    .X(net3586));
 sky130_fd_sc_hs__buf_1 place3613 (.A(net3612),
    .X(net3613));
 sky130_fd_sc_hs__buf_1 place3621 (.A(_02204_),
    .X(net3621));
 sky130_fd_sc_hs__buf_1 place3623 (.A(net3622),
    .X(net3623));
 sky130_fd_sc_hs__buf_1 place3627 (.A(net3626),
    .X(net3627));
 sky130_fd_sc_hs__buf_1 place3636 (.A(_02108_),
    .X(net3636));
 sky130_fd_sc_hs__buf_1 place3650 (.A(_02048_),
    .X(net3650));
 sky130_fd_sc_hs__buf_1 place3658 (.A(net3657),
    .X(net3658));
 sky130_fd_sc_hs__buf_1 place3675 (.A(_00589_),
    .X(net3675));
 sky130_fd_sc_hs__buf_1 place3676 (.A(\u_window_buffer.write_ptr[9] ),
    .X(net3676));
 sky130_fd_sc_hs__buf_1 place3677 (.A(\u_window_buffer.write_ptr[9] ),
    .X(net3677));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__inv_16 clkload0 (.A(clknet_2_1__leaf_clk));
 sky130_fd_sc_hs__clkinv_16 clkload1 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hs__inv_16 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hs__clkbuf_16 clkload3 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hs__clkinv_1 clkload4 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hs__clkbuf_16 clkload5 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hs__clkinv_1 clkload6 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hs__clkbuf_16 clkload7 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hs__clkinv_1 clkload8 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hs__clkinv_2 clkload9 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hs__clkbuf_16 clkload10 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hs__clkbuf_8 clkload11 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hs__clkinv_4 clkload12 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hs__clkinv_1 clkload13 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hs__clkbuf_16 clkload14 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hs__clkinv_4 clkload15 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hs__clkinv_2 clkload16 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hs__clkbuf_16 clkload17 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hs__clkinv_2 clkload18 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hs__clkinv_2 clkload19 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hs__clkinv_2 clkload20 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hs__clkinv_1 clkload21 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hs__clkinv_4 clkload22 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hs__clkinv_2 clkload23 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hs__clkinv_2 clkload24 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hs__clkbuf_16 clkload25 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hs__clkinv_2 clkload26 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hs__clkinv_2 clkload27 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hs__clkinv_2 clkload28 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hs__clkbuf_16 clkload29 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hs__clkinv_1 clkload30 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hs__clkinv_4 clkload31 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hs__clkinv_2 clkload32 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hs__clkinv_1 clkload33 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hs__clkbuf_2 clkload34 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hs__clkinv_1 clkload35 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hs__nand2_8 clone3786 (.A(net3787),
    .B(net2966),
    .Y(net3786));
 sky130_fd_sc_hs__buf_8 rebuffer3787 (.A(_01962_),
    .X(net3787));
 sky130_fd_sc_hs__clkbuf_16 rebuffer3788 (.A(_04775_),
    .X(net3788));
 sky130_fd_sc_hs__buf_4 rebuffer3789 (.A(_00136_),
    .X(net3789));
 sky130_fd_sc_hs__buf_1 rebuffer3790 (.A(_00883_),
    .X(net3790));
 sky130_fd_sc_hs__buf_1 rebuffer3791 (.A(_00828_),
    .X(net3791));
 sky130_fd_sc_hs__buf_1 rebuffer3792 (.A(_01216_),
    .X(net3792));
 sky130_fd_sc_hs__buf_1 rebuffer3793 (.A(_01749_),
    .X(net3793));
 sky130_fd_sc_hs__buf_2 rebuffer3794 (.A(_01901_),
    .X(net3794));
 sky130_fd_sc_hs__buf_1 rebuffer3795 (.A(_01455_),
    .X(net3795));
 sky130_fd_sc_hs__buf_1 rebuffer3796 (.A(net3805),
    .X(net3796));
 sky130_fd_sc_hs__buf_1 rebuffer3797 (.A(_01743_),
    .X(net3797));
 sky130_fd_sc_hs__buf_1 rebuffer3798 (.A(_01577_),
    .X(net3798));
 sky130_fd_sc_hs__buf_1 rebuffer3799 (.A(_01715_),
    .X(net3799));
 sky130_fd_sc_hs__buf_1 rebuffer3800 (.A(_01552_),
    .X(net3800));
 sky130_fd_sc_hs__buf_8 rebuffer3801 (.A(_00987_),
    .X(net3801));
 sky130_fd_sc_hs__buf_1 rebuffer3802 (.A(_01264_),
    .X(net3802));
 sky130_fd_sc_hs__buf_1 rebuffer3803 (.A(_01880_),
    .X(net3803));
 sky130_fd_sc_hs__buf_1 rebuffer3804 (.A(_01657_),
    .X(net3804));
 sky130_fd_sc_hs__buf_2 rebuffer3805 (.A(_01743_),
    .X(net3805));
 sky130_fd_sc_hs__buf_1 rebuffer3806 (.A(_01306_),
    .X(net3806));
 sky130_fd_sc_hs__buf_1 rebuffer3832 (.A(_01641_),
    .X(net3832));
 sky130_fd_sc_hs__buf_1 rebuffer3833 (.A(_01355_),
    .X(net3833));
 sky130_fd_sc_hs__buf_1 rebuffer3834 (.A(_01839_),
    .X(net3834));
 sky130_fd_sc_hs__buf_1 rebuffer3835 (.A(_01839_),
    .X(net3835));
 sky130_fd_sc_hs__buf_1 rebuffer3836 (.A(_01839_),
    .X(net3836));
 sky130_fd_sc_hs__buf_1 rebuffer3837 (.A(_01820_),
    .X(net3837));
 sky130_fd_sc_hs__buf_1 rebuffer3838 (.A(_01164_),
    .X(net3838));
 sky130_fd_sc_hs__buf_1 rebuffer3839 (.A(_01425_),
    .X(net3839));
 sky130_fd_sc_hs__buf_1 rebuffer3840 (.A(_01425_),
    .X(net3840));
 sky130_fd_sc_hs__buf_1 rebuffer3841 (.A(_01361_),
    .X(net3841));
 sky130_fd_sc_hs__buf_1 rebuffer4860 (.A(_04438_),
    .X(net4860));
 sky130_fd_sc_hs__buf_1 rebuffer4861 (.A(_04438_),
    .X(net4861));
 sky130_fd_sc_hs__buf_1 rebuffer4862 (.A(_01216_),
    .X(net4862));
 sky130_fd_sc_hs__buf_1 rebuffer4863 (.A(_01373_),
    .X(net4863));
 sky130_fd_sc_hs__buf_2 rebuffer4864 (.A(_01228_),
    .X(net4864));
 sky130_fd_sc_hs__buf_1 rebuffer4865 (.A(_01216_),
    .X(net4865));
 sky130_fd_sc_hs__buf_1 rebuffer4866 (.A(_01489_),
    .X(net4866));
 sky130_fd_sc_hs__buf_1 rebuffer4867 (.A(_01878_),
    .X(net4867));
 sky130_fd_sc_hs__buf_1 rebuffer4868 (.A(_01160_),
    .X(net4868));
 sky130_fd_sc_hs__buf_1 rebuffer4869 (.A(_00931_),
    .X(net4869));
 sky130_fd_sc_hs__buf_1 rebuffer4870 (.A(_00931_),
    .X(net4870));
 sky130_fd_sc_hs__buf_1 rebuffer4871 (.A(_01633_),
    .X(net4871));
 sky130_fd_sc_hs__buf_1 rebuffer4872 (.A(_01369_),
    .X(net4872));
 sky130_fd_sc_hs__buf_1 rebuffer4873 (.A(_01934_),
    .X(net4873));
 sky130_fd_sc_hs__buf_1 rebuffer4874 (.A(_00894_),
    .X(net4874));
 sky130_fd_sc_hs__buf_2 rebuffer4875 (.A(_00728_),
    .X(net4875));
 sky130_fd_sc_hs__buf_1 rebuffer4876 (.A(net4875),
    .X(net4876));
 sky130_fd_sc_hs__buf_2 rebuffer4877 (.A(_00977_),
    .X(net4877));
 sky130_fd_sc_hs__buf_1 rebuffer4888 (.A(_04015_),
    .X(net4888));
 sky130_fd_sc_hs__buf_1 rebuffer4889 (.A(_04782_),
    .X(net4889));
 sky130_fd_sc_hs__buf_1 rebuffer4890 (.A(_04617_),
    .X(net4890));
 sky130_fd_sc_hs__buf_1 rebuffer4891 (.A(_04013_),
    .X(net4891));
 sky130_fd_sc_hs__buf_1 rebuffer4892 (.A(_01765_),
    .X(net4892));
 sky130_fd_sc_hs__buf_1 rebuffer4893 (.A(_01901_),
    .X(net4893));
 sky130_fd_sc_hs__buf_1 rebuffer4894 (.A(_01960_),
    .X(net4894));
 sky130_fd_sc_hs__buf_1 rebuffer4895 (.A(_01233_),
    .X(net4895));
 sky130_fd_sc_hs__buf_1 rebuffer4896 (.A(_01600_),
    .X(net4896));
 sky130_fd_sc_hs__buf_1 rebuffer4897 (.A(_01353_),
    .X(net4897));
 sky130_fd_sc_hs__buf_1 rebuffer4898 (.A(_01892_),
    .X(net4898));
 sky130_fd_sc_hs__buf_1 rebuffer4899 (.A(_04042_),
    .X(net4899));
 sky130_fd_sc_hs__buf_2 rebuffer4900 (.A(_04587_),
    .X(net4900));
 sky130_fd_sc_hs__buf_1 rebuffer4901 (.A(_04587_),
    .X(net4901));
 sky130_fd_sc_hs__buf_1 rebuffer4902 (.A(_01798_),
    .X(net4902));
 sky130_fd_sc_hs__buf_2 rebuffer4903 (.A(net1848),
    .X(net4903));
 sky130_fd_sc_hs__buf_1 rebuffer4904 (.A(_01670_),
    .X(net4904));
 sky130_fd_sc_hs__buf_1 rebuffer4905 (.A(_00853_),
    .X(net4905));
 sky130_fd_sc_hs__buf_1 rebuffer4906 (.A(_04561_),
    .X(net4906));
 sky130_fd_sc_hs__buf_1 rebuffer4907 (.A(_01306_),
    .X(net4907));
 sky130_fd_sc_hs__buf_1 rebuffer4908 (.A(_01504_),
    .X(net4908));
 sky130_fd_sc_hs__buf_1 rebuffer4918 (.A(_01545_),
    .X(net4918));
 sky130_fd_sc_hs__buf_1 rebuffer4919 (.A(_01522_),
    .X(net4919));
 sky130_fd_sc_hs__buf_1 rebuffer4920 (.A(_01504_),
    .X(net4920));
 sky130_fd_sc_hs__buf_1 rebuffer4921 (.A(_00932_),
    .X(net4921));
 sky130_fd_sc_hs__buf_1 rebuffer4922 (.A(_01056_),
    .X(net4922));
 sky130_fd_sc_hs__buf_1 rebuffer4924 (.A(_01311_),
    .X(net4924));
 sky130_fd_sc_hs__buf_1 rebuffer4925 (.A(_00729_),
    .X(net4925));
 sky130_fd_sc_hs__buf_1 rebuffer4926 (.A(_00828_),
    .X(net4926));
 sky130_fd_sc_hs__buf_1 rebuffer4927 (.A(_01490_),
    .X(net4927));
 sky130_fd_sc_hs__buf_1 rebuffer4928 (.A(_01956_),
    .X(net4928));
 sky130_fd_sc_hs__buf_1 rebuffer4929 (.A(_01635_),
    .X(net4929));
 sky130_fd_sc_hs__buf_1 rebuffer4930 (.A(_01635_),
    .X(net4930));
 sky130_fd_sc_hs__buf_1 rebuffer4931 (.A(_01866_),
    .X(net4931));
 sky130_fd_sc_hs__bufbuf_8 rebuffer4932 (.A(_01738_),
    .X(net4932));
 sky130_fd_sc_hs__buf_1 rebuffer4933 (.A(_00906_),
    .X(net4933));
 sky130_fd_sc_hs__buf_8 rebuffer4934 (.A(net3786),
    .X(net4934));
 sky130_fd_sc_hs__buf_16 clone4962 (.A(net4967),
    .X(net4962));
 sky130_fd_sc_hs__buf_16 rebuffer4967 (.A(net1845),
    .X(net4967));
 sky130_fd_sc_hs__buf_8 clone4972 (.A(_04775_),
    .X(net4972));
 sky130_fd_sc_hs__buf_16 clone4973 (.A(net4967),
    .X(net4973));
 sky130_fd_sc_hs__buf_16 clone4974 (.A(net4975),
    .X(net4974));
 sky130_fd_sc_hs__buf_8 rebuffer4975 (.A(_04792_),
    .X(net4975));
 sky130_fd_sc_hs__buf_8 rebuffer5040 (.A(net1844),
    .X(net5040));
 sky130_fd_sc_hs__clkbuf_2 rebuffer5041 (.A(net1844),
    .X(net5041));
 sky130_fd_sc_hs__buf_1 rebuffer5042 (.A(_04879_),
    .X(net5042));
 sky130_fd_sc_hs__buf_1 rebuffer5043 (.A(_05517_),
    .X(net5043));
 sky130_fd_sc_hs__buf_8 clone5044 (.A(_05722_),
    .X(net5044));
 sky130_fd_sc_hs__buf_1 rebuffer5045 (.A(_05211_),
    .X(net5045));
 sky130_fd_sc_hs__buf_1 rebuffer5046 (.A(_05211_),
    .X(net5046));
 sky130_fd_sc_hs__bufbuf_8 rebuffer5047 (.A(_05171_),
    .X(net5047));
 sky130_fd_sc_hs__buf_1 rebuffer5048 (.A(_05143_),
    .X(net5048));
 sky130_fd_sc_hs__buf_1 rebuffer5049 (.A(_05431_),
    .X(net5049));
 sky130_fd_sc_hs__buf_2 rebuffer5050 (.A(_05431_),
    .X(net5050));
 sky130_fd_sc_hs__clkbuf_2 rebuffer5051 (.A(_05360_),
    .X(net5051));
 sky130_fd_sc_hs__buf_1 rebuffer5052 (.A(_05217_),
    .X(net5052));
 sky130_fd_sc_hs__buf_1 rebuffer5053 (.A(_05041_),
    .X(net5053));
 sky130_fd_sc_hs__buf_1 rebuffer5054 (.A(_05427_),
    .X(net5054));
 sky130_fd_sc_hs__buf_1 rebuffer5055 (.A(_05674_),
    .X(net5055));
 sky130_fd_sc_hs__buf_1 rebuffer5056 (.A(_04901_),
    .X(net5056));
 sky130_fd_sc_hs__buf_1 rebuffer5057 (.A(_04838_),
    .X(net5057));
 sky130_fd_sc_hs__buf_2 rebuffer5058 (.A(_05247_),
    .X(net5058));
 sky130_fd_sc_hs__buf_1 rebuffer5059 (.A(_05273_),
    .X(net5059));
 sky130_fd_sc_hs__buf_1 rebuffer5060 (.A(_05039_),
    .X(net5060));
 sky130_fd_sc_hs__buf_1 rebuffer5061 (.A(_04827_),
    .X(net5061));
 sky130_fd_sc_hs__buf_1 rebuffer5062 (.A(_05605_),
    .X(net5062));
 sky130_fd_sc_hs__buf_1 rebuffer5063 (.A(_04885_),
    .X(net5063));
 sky130_fd_sc_hs__buf_1 rebuffer5064 (.A(_05100_),
    .X(net5064));
 sky130_fd_sc_hs__buf_1 rebuffer5066 (.A(_05096_),
    .X(net5066));
 sky130_fd_sc_hs__buf_1 rebuffer5067 (.A(_05153_),
    .X(net5067));
 sky130_fd_sc_hs__buf_1 rebuffer5068 (.A(_05427_),
    .X(net5068));
 sky130_fd_sc_hs__buf_1 rebuffer5069 (.A(_05035_),
    .X(net5069));
 sky130_fd_sc_hs__buf_1 rebuffer5070 (.A(_05029_),
    .X(net5070));
 sky130_fd_sc_hs__buf_1 rebuffer5071 (.A(_05721_),
    .X(net5071));
 sky130_fd_sc_hs__buf_1 rebuffer5072 (.A(_05355_),
    .X(net5072));
 sky130_fd_sc_hs__buf_1 rebuffer5073 (.A(_05312_),
    .X(net5073));
 sky130_fd_sc_hs__buf_2 rebuffer5074 (.A(_05480_),
    .X(net5074));
 sky130_fd_sc_hs__buf_1 rebuffer5075 (.A(\u_window_buffer.write_ptr[0] ),
    .X(net5075));
 sky130_fd_sc_hs__buf_1 rebuffer5076 (.A(_04827_),
    .X(net5076));
 sky130_fd_sc_hs__buf_1 rebuffer5077 (.A(_05305_),
    .X(net5077));
 sky130_fd_sc_hs__buf_1 rebuffer5078 (.A(_05029_),
    .X(net5078));
 sky130_fd_sc_hs__buf_1 rebuffer5079 (.A(_05168_),
    .X(net5079));
 sky130_fd_sc_hs__buf_1 rebuffer5080 (.A(_05365_),
    .X(net5080));
 sky130_fd_sc_hs__buf_1 rebuffer5081 (.A(_04939_),
    .X(net5081));
 sky130_fd_sc_hs__buf_1 rebuffer5082 (.A(_05274_),
    .X(net5082));
 sky130_fd_sc_hs__buf_1 rebuffer5083 (.A(net2031),
    .X(net5083));
 sky130_fd_sc_hs__buf_8 rebuffer5084 (.A(_05697_),
    .X(net5084));
 sky130_fd_sc_hs__buf_1 rebuffer5085 (.A(_05128_),
    .X(net5085));
 sky130_fd_sc_hs__buf_1 rebuffer5086 (.A(_04826_),
    .X(net5086));
 sky130_fd_sc_hs__buf_1 rebuffer5087 (.A(_05506_),
    .X(net5087));
 sky130_fd_sc_hs__buf_1 rebuffer5088 (.A(_05512_),
    .X(net5088));
 sky130_fd_sc_hs__buf_1 rebuffer5090 (.A(_05004_),
    .X(net5090));
 sky130_fd_sc_hs__buf_1 rebuffer5091 (.A(_05585_),
    .X(net5091));
 sky130_fd_sc_hs__buf_1 rebuffer5092 (.A(_05031_),
    .X(net5092));
 sky130_fd_sc_hs__buf_1 rebuffer5093 (.A(net2191),
    .X(net5093));
 sky130_fd_sc_hs__buf_1 rebuffer5094 (.A(net2191),
    .X(net5094));
 sky130_fd_sc_hs__buf_1 rebuffer5095 (.A(_05486_),
    .X(net5095));
 sky130_fd_sc_hs__buf_1 rebuffer5097 (.A(_05099_),
    .X(net5097));
 sky130_fd_sc_hs__buf_1 rebuffer5098 (.A(_05642_),
    .X(net5098));
 sky130_fd_sc_hs__buf_1 rebuffer5099 (.A(_05290_),
    .X(net5099));
 sky130_fd_sc_hs__buf_1 rebuffer5100 (.A(_05580_),
    .X(net5100));
 sky130_fd_sc_hs__buf_1 rebuffer5101 (.A(_05346_),
    .X(net5101));
 sky130_fd_sc_hs__buf_1 rebuffer5102 (.A(_05262_),
    .X(net5102));
 sky130_fd_sc_hs__buf_1 rebuffer5103 (.A(net2471),
    .X(net5103));
 sky130_fd_sc_hs__buf_1 rebuffer5104 (.A(_05271_),
    .X(net5104));
 sky130_fd_sc_hs__buf_16 clone5105 (.A(net5106),
    .X(net5105));
 sky130_fd_sc_hs__buf_8 rebuffer5106 (.A(_05708_),
    .X(net5106));
 sky130_fd_sc_hs__buf_1 rebuffer5108 (.A(_03263_),
    .X(net5108));
 sky130_fd_sc_hs__buf_1 rebuffer5109 (.A(_03582_),
    .X(net5109));
 sky130_fd_sc_hs__buf_1 rebuffer5110 (.A(_03120_),
    .X(net5110));
 sky130_fd_sc_hs__buf_1 rebuffer5111 (.A(net5110),
    .X(net5111));
 sky130_fd_sc_hs__buf_1 rebuffer5112 (.A(_03120_),
    .X(net5112));
 sky130_fd_sc_hs__buf_1 rebuffer5113 (.A(_03182_),
    .X(net5113));
 sky130_fd_sc_hs__buf_1 rebuffer5114 (.A(_03182_),
    .X(net5114));
 sky130_fd_sc_hs__buf_1 rebuffer5115 (.A(_03213_),
    .X(net5115));
 sky130_fd_sc_hs__buf_2 rebuffer5116 (.A(_03064_),
    .X(net5116));
 sky130_fd_sc_hs__buf_1 rebuffer5117 (.A(_03064_),
    .X(net5117));
 sky130_fd_sc_hs__buf_1 rebuffer5118 (.A(_03493_),
    .X(net5118));
 sky130_fd_sc_hs__buf_1 rebuffer5119 (.A(_03593_),
    .X(net5119));
 sky130_fd_sc_hs__buf_1 rebuffer5120 (.A(_03493_),
    .X(net5120));
 sky130_fd_sc_hs__buf_1 rebuffer5121 (.A(_03006_),
    .X(net5121));
 sky130_fd_sc_hs__buf_2 rebuffer5122 (.A(_03177_),
    .X(net5122));
 sky130_fd_sc_hs__buf_1 rebuffer5123 (.A(_02878_),
    .X(net5123));
 sky130_fd_sc_hs__buf_1 rebuffer5124 (.A(_02958_),
    .X(net5124));
 sky130_fd_sc_hs__buf_1 rebuffer5125 (.A(_03031_),
    .X(net5125));
 sky130_fd_sc_hs__buf_2 rebuffer5126 (.A(_03582_),
    .X(net5126));
 sky130_fd_sc_hs__buf_1 rebuffer5127 (.A(_02941_),
    .X(net5127));
 sky130_fd_sc_hs__buf_1 rebuffer5128 (.A(_03529_),
    .X(net5128));
 sky130_fd_sc_hs__buf_1 rebuffer5129 (.A(_03009_),
    .X(net5129));
 sky130_fd_sc_hs__buf_1 rebuffer5130 (.A(_03408_),
    .X(net5130));
 sky130_fd_sc_hs__buf_1 rebuffer5131 (.A(_03554_),
    .X(net5131));
 sky130_fd_sc_hs__buf_1 rebuffer5132 (.A(_03017_),
    .X(net5132));
 sky130_fd_sc_hs__buf_1 rebuffer5133 (.A(_03526_),
    .X(net5133));
 sky130_fd_sc_hs__buf_1 rebuffer5134 (.A(_03181_),
    .X(net5134));
 sky130_fd_sc_hs__buf_2 rebuffer5135 (.A(_03658_),
    .X(net5135));
 sky130_fd_sc_hs__buf_1 rebuffer5136 (.A(_03364_),
    .X(net5136));
 sky130_fd_sc_hs__buf_2 rebuffer5137 (.A(_03215_),
    .X(net5137));
 sky130_fd_sc_hs__buf_2 rebuffer5138 (.A(_03245_),
    .X(net5138));
 sky130_fd_sc_hs__buf_1 rebuffer5139 (.A(_03366_),
    .X(net5139));
 sky130_fd_sc_hs__buf_2 rebuffer5140 (.A(_03366_),
    .X(net5140));
 sky130_fd_sc_hs__buf_1 rebuffer5141 (.A(_03112_),
    .X(net5141));
 sky130_fd_sc_hs__buf_1 rebuffer5143 (.A(_03097_),
    .X(net5143));
 sky130_fd_sc_hs__buf_1 rebuffer5144 (.A(_02944_),
    .X(net5144));
 sky130_fd_sc_hs__buf_1 rebuffer5165 (.A(_03396_),
    .X(net5165));
 sky130_fd_sc_hs__buf_1 rebuffer5166 (.A(_03348_),
    .X(net5166));
 sky130_fd_sc_hs__buf_2 rebuffer5167 (.A(_03213_),
    .X(net5167));
 sky130_fd_sc_hs__buf_1 rebuffer5168 (.A(_02996_),
    .X(net5168));
 sky130_fd_sc_hs__buf_1 rebuffer5169 (.A(_03022_),
    .X(net5169));
 sky130_fd_sc_hs__buf_1 rebuffer5170 (.A(_02981_),
    .X(net5170));
 sky130_fd_sc_hs__buf_1 rebuffer5171 (.A(_03227_),
    .X(net5171));
 sky130_fd_sc_hs__buf_1 rebuffer5172 (.A(_03230_),
    .X(net5172));
 sky130_fd_sc_hs__buf_2 rebuffer5173 (.A(_03159_),
    .X(net5173));
 sky130_fd_sc_hs__buf_1 rebuffer5174 (.A(net3749),
    .X(net5174));
 sky130_fd_sc_hs__buf_1 rebuffer5175 (.A(_03308_),
    .X(net5175));
 sky130_fd_sc_hs__buf_1 rebuffer5176 (.A(net3301),
    .X(net5176));
 sky130_fd_sc_hs__buf_4 rebuffer5177 (.A(_03339_),
    .X(net5177));
 sky130_fd_sc_hs__buf_1 rebuffer5178 (.A(_03229_),
    .X(net5178));
 sky130_fd_sc_hs__buf_1 rebuffer5179 (.A(_03169_),
    .X(net5179));
 sky130_fd_sc_hs__buf_1 rebuffer5180 (.A(_03161_),
    .X(net5180));
 sky130_fd_sc_hs__buf_4 rebuffer5181 (.A(_03274_),
    .X(net5181));
 sky130_fd_sc_hs__buf_1 rebuffer5182 (.A(_03204_),
    .X(net5182));
 sky130_fd_sc_hs__buf_1 rebuffer5183 (.A(_00220_),
    .X(net5183));
 sky130_fd_sc_hs__buf_1 rebuffer5191 (.A(_03640_),
    .X(net5191));
 sky130_fd_sc_hs__buf_1 rebuffer5192 (.A(_03246_),
    .X(net5192));
 sky130_fd_sc_hs__buf_1 rebuffer5193 (.A(_03029_),
    .X(net5193));
 sky130_fd_sc_hs__buf_1 rebuffer5194 (.A(_03029_),
    .X(net5194));
 sky130_fd_sc_hs__buf_1 rebuffer5195 (.A(net3301),
    .X(net5195));
 sky130_fd_sc_hs__buf_1 rebuffer5196 (.A(_03335_),
    .X(net5196));
 sky130_fd_sc_hs__buf_1 rebuffer5199 (.A(_05719_),
    .X(net5199));
endmodule
