module FFT #(
    parameter NFFT = 512
) (
    input  logic clk,
    input  logic rst_n,
);
    
endmodule