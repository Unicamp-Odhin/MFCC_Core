`timescale 1ns/1ps

module FFT #(
    parameter NFFT = 512
) (
    input  logic clk,
    input  logic rst_n,
);
    
endmodule