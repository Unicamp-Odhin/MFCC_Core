`timescale 1ns/1ps

module DCT #(
    parameter NUM_CEPS = 12
) (
    input  logic clk,
    input  logic rst_n,
);

logic signed [15:0] cos_table [40][12] = '{
    '{ 32767, 32742, 32666, 32540, 32364, 32138, 31862, 31537, 31164, 30742, 30273, 29758 },
    '{ 32767, 32540, 31862, 30742, 29196, 27245, 24916, 22242, 19260, 16011, 12539, 8894 },
    '{ 32767, 32138, 30273, 27245, 23170, 18204, 12539, 6392, 0, -6392, -12539, -18204 },
    '{ 32767, 31537, 27939, 22242, 14876, 6392, -2570, -11341, -19260, -25733, -30273, -32540 },
    '{ 32767, 30742, 24916, 16011, 5126, -6392, -17121, -25733, -31164, -32742, -30273, -24062 },
    '{ 32767, 29758, 21281, 8894, -5126, -18204, -27939, -32540, -31164, -24062, -12539, 1286 },
    '{ 32767, 28589, 17121, 1286, -14876, -27245, -32666, -29758, -19260, -3851, 12539, 25733 },
    '{ 32767, 27245, 12539, -6392, -23170, -32138, -30273, -18204, 0, 18204, 30273, 32138 },
    '{ 32767, 25733, 7649, -13718, -29196, -32138, -21281, -1286, 19260, 31537, 30273, 16011 },
    '{ 32767, 24062, 2570, -20286, -32364, -27245, -7649, 16011, 31164, 29758, 12539, -11341 },
    '{ 32767, 22242, -2570, -25733, -32364, -18204, 7649, 28589, 31164, 13718, -12539, -30742 },
    '{ 32767, 20286, -7649, -29758, -29196, -6392, 21281, 32742, 19260, -8894, -30273, -28589 },
    '{ 32767, 18204, -12539, -32138, -23170, 6392, 30273, 27245, 0, -27245, -30273, -6392 },
    '{ 32767, 16011, -17121, -32742, -14876, 18204, 32666, 13718, -19260, -32540, -12539, 20286 },
    '{ 32767, 13718, -21281, -31537, -5126, 27245, 27939, -3851, -31164, -22242, 12539, 32742 },
    '{ 32767, 11341, -24916, -28589, 5126, 32138, 17121, -20286, -31164, -1286, 30273, 22242 },
    '{ 32767, 8894, -27939, -24062, 14876, 32138, 2570, -30742, -19260, 20286, 30273, -3851 },
    '{ 32767, 6392, -30273, -18204, 23170, 27245, -12539, -32138, 0, 32138, 12539, -27245 },
    '{ 32767, 3851, -31862, -11341, 29196, 18204, -24916, -24062, 19260, 28589, -12539, -31537 },
    '{ 32767, 1286, -32666, -3851, 32364, 6392, -31862, -8894, 31164, 11341, -30273, -13718 },
    '{ 32767, -1286, -32666, 3851, 32364, -6392, -31862, 8894, 31164, -11341, -30273, 13718 },
    '{ 32767, -3851, -31862, 11341, 29196, -18204, -24916, 24062, 19260, -28589, -12539, 31537 },
    '{ 32767, -6392, -30273, 18204, 23170, -27245, -12539, 32138, 0, -32138, 12539, 27245 },
    '{ 32767, -8894, -27939, 24062, 14876, -32138, 2570, 30742, -19260, -20286, 30273, 3851 },
    '{ 32767, -11341, -24916, 28589, 5126, -32138, 17121, 20286, -31164, 1286, 30273, -22242 },
    '{ 32767, -13718, -21281, 31537, -5126, -27245, 27939, 3851, -31164, 22242, 12539, -32742 },
    '{ 32767, -16011, -17121, 32742, -14876, -18204, 32666, -13718, -19260, 32540, -12539, -20286 },
    '{ 32767, -18204, -12539, 32138, -23170, -6392, 30273, -27245, 0, 27245, -30273, 6392 },
    '{ 32767, -20286, -7649, 29758, -29196, 6392, 21281, -32742, 19260, 8894, -30273, 28589 },
    '{ 32767, -22242, -2570, 25733, -32364, 18204, 7649, -28589, 31164, -13718, -12539, 30742 },
    '{ 32767, -24062, 2570, 20286, -32364, 27245, -7649, -16011, 31164, -29758, 12539, 11341 },
    '{ 32767, -25733, 7649, 13718, -29196, 32138, -21281, 1286, 19260, -31537, 30273, -16011 },
    '{ 32767, -27245, 12539, 6392, -23170, 32138, -30273, 18204, 0, -18204, 30273, -32138 },
    '{ 32767, -28589, 17121, -1286, -14876, 27245, -32666, 29758, -19260, 3851, 12539, -25733 },
    '{ 32767, -29758, 21281, -8894, -5126, 18204, -27939, 32540, -31164, 24062, -12539, -1286 },
    '{ 32767, -30742, 24916, -16011, 5126, 6392, -17121, 25733, -31164, 32742, -30273, 24062 },
    '{ 32767, -31537, 27939, -22242, 14876, -6392, -2570, 11341, -19260, 25733, -30273, 32540 },
    '{ 32767, -32138, 30273, -27245, 23170, -18204, 12539, -6392, 0, 6392, -12539, 18204 },
    '{ 32767, -32540, 31862, -30742, 29196, -27245, 24916, -22242, 19260, -16011, 12539, -8894 },
    '{ 32767, -32742, 32666, -32540, 32364, -32138, 31862, -31537, 31164, -30742, 30273, -29758 }
};

endmodule