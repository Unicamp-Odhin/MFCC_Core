module MFCC_Core (auto_restart_i,
    clk,
    mfcc_done_o,
    pcm_ready_i,
    rst_n,
    start_i,
    mfcc_data_o,
    pcm_in);
 input auto_restart_i;
 input clk;
 output mfcc_done_o;
 input pcm_ready_i;
 input rst_n;
 input start_i;
 output [207:0] mfcc_data_o;
 input [15:0] pcm_in;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire net3054;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire net3053;
 wire net3052;
 wire net3058;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire net3051;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire net3050;
 wire net3049;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire net3047;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire net3046;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire net3045;
 wire _00958_;
 wire net3043;
 wire _00960_;
 wire net3042;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire net3041;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire net3040;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire net3044;
 wire net3039;
 wire _01012_;
 wire net3038;
 wire _01014_;
 wire _01015_;
 wire net3037;
 wire _01017_;
 wire net3036;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire net3035;
 wire _01024_;
 wire _01025_;
 wire net3034;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire net3033;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire net3032;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire net3031;
 wire net3030;
 wire _01080_;
 wire _01081_;
 wire net3029;
 wire net3028;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire net3048;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire net3026;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire net3025;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire net3024;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire net3023;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire net3022;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire net3021;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire net3020;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire net3018;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire net3017;
 wire net3016;
 wire _02511_;
 wire net3019;
 wire _02513_;
 wire _02514_;
 wire net3015;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire net3027;
 wire net3012;
 wire _02527_;
 wire net3011;
 wire net3010;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire net3009;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire net3008;
 wire net3007;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire net3005;
 wire _02603_;
 wire _02604_;
 wire net3003;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire net3001;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire net3002;
 wire _02654_;
 wire net3004;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire net3000;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire net2999;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire net2998;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire net2997;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire net2996;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire net2995;
 wire _02853_;
 wire _02854_;
 wire net2994;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire net2993;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire net2992;
 wire _02866_;
 wire _02867_;
 wire net2991;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire net2990;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire net3006;
 wire _02879_;
 wire _02880_;
 wire net2988;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire net2987;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire net2986;
 wire _02899_;
 wire net2985;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire net2984;
 wire net2983;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire net2982;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire net2981;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire net2980;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire net2979;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire net2978;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire net2989;
 wire net2976;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire net2977;
 wire _03162_;
 wire net2975;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire net2974;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire net2973;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire net2972;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire net2971;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire net2970;
 wire _04153_;
 wire net2969;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire net2968;
 wire _04165_;
 wire net2966;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire net2965;
 wire net2964;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire net2962;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire net2961;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire net2960;
 wire net2959;
 wire _04333_;
 wire net2956;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire net2955;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire net2954;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire net2953;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire net2952;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire net2951;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire net2957;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire net2950;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire net2949;
 wire _05374_;
 wire _05375_;
 wire net2946;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire net2944;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire net2942;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire net2941;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire net2940;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire net2939;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire net2938;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire net2937;
 wire net2936;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire net2934;
 wire net2933;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire net2932;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire net2930;
 wire _06484_;
 wire net2929;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire net2931;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire net3055;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire \mel_ptr[0] ;
 wire \mel_ptr[1] ;
 wire net213;
 wire \tx_fifo.read_ptr[0] ;
 wire \tx_fifo.read_ptr[1] ;
 wire \tx_fifo.write_ptr[0] ;
 wire \tx_fifo.write_ptr[1] ;
 wire \u_dct.k_ptr[0] ;
 wire \u_dct.k_ptr[1] ;
 wire \u_dct.n_ptr[0] ;
 wire \u_dct.n_ptr[1] ;
 wire \u_fft.power_ptr[0] ;
 wire \u_fft.power_ptr[1] ;
 wire \u_fft.sched[30] ;
 wire \u_fft.sched[31] ;
 wire \u_fft.sched[32] ;
 wire \u_fft.sched[33] ;
 wire \u_fft.sched[34] ;
 wire \u_fft.sched[35] ;
 wire \u_fft.sched[36] ;
 wire \u_fft.sched[37] ;
 wire \u_fft.sched[38] ;
 wire \u_fft.sched[40] ;
 wire \u_fft.sched[41] ;
 wire \u_fft.sched[42] ;
 wire \u_fft.sched[45] ;
 wire \u_fft.sched[46] ;
 wire \u_fft.sched[47] ;
 wire \u_fft.sched[48] ;
 wire \u_fft.sched[49] ;
 wire \u_fft.sched[50] ;
 wire \u_fft.sched[51] ;
 wire \u_fft.sched[52] ;
 wire \u_fft.sched[53] ;
 wire \u_fft.sched[54] ;
 wire \u_fft.sched[55] ;
 wire \u_fft.sched[56] ;
 wire \u_fft.sched[57] ;
 wire \u_fft.sched[58] ;
 wire \u_fft.sched[59] ;
 wire \u_fft.sched[60] ;
 wire \u_fft.sched[61] ;
 wire \u_fft.sched[62] ;
 wire \u_fft.sched[63] ;
 wire \u_fft.sched[64] ;
 wire \u_hamming_window.calc_pointer[0] ;
 wire \u_hamming_window.calc_pointer[1] ;
 wire \u_hamming_window.done ;
 wire \u_hamming_window.frame_ptr[0] ;
 wire \u_hamming_window.frame_ptr[1] ;
 wire \u_mel.k[0] ;
 wire \u_mel.k[1] ;
 wire \u_mel.k_next[0] ;
 wire \u_window_buffer.internal_read_ptr[10] ;
 wire \u_window_buffer.internal_read_ptr[11] ;
 wire \u_window_buffer.internal_read_ptr[12] ;
 wire \u_window_buffer.internal_read_ptr[13] ;
 wire \u_window_buffer.internal_read_ptr[14] ;
 wire \u_window_buffer.internal_read_ptr[15] ;
 wire \u_window_buffer.internal_read_ptr[16] ;
 wire \u_window_buffer.internal_read_ptr[17] ;
 wire \u_window_buffer.internal_read_ptr[18] ;
 wire \u_window_buffer.internal_read_ptr[19] ;
 wire \u_window_buffer.internal_read_ptr[1] ;
 wire \u_window_buffer.internal_read_ptr[20] ;
 wire \u_window_buffer.internal_read_ptr[21] ;
 wire \u_window_buffer.internal_read_ptr[22] ;
 wire \u_window_buffer.internal_read_ptr[23] ;
 wire \u_window_buffer.internal_read_ptr[24] ;
 wire \u_window_buffer.internal_read_ptr[25] ;
 wire \u_window_buffer.internal_read_ptr[26] ;
 wire \u_window_buffer.internal_read_ptr[27] ;
 wire \u_window_buffer.internal_read_ptr[28] ;
 wire \u_window_buffer.internal_read_ptr[29] ;
 wire \u_window_buffer.internal_read_ptr[2] ;
 wire \u_window_buffer.internal_read_ptr[30] ;
 wire \u_window_buffer.internal_read_ptr[3] ;
 wire \u_window_buffer.internal_read_ptr[4] ;
 wire \u_window_buffer.internal_read_ptr[5] ;
 wire \u_window_buffer.internal_read_ptr[6] ;
 wire \u_window_buffer.internal_read_ptr[7] ;
 wire \u_window_buffer.internal_read_ptr[8] ;
 wire \u_window_buffer.internal_read_ptr[9] ;
 wire \u_window_buffer.move_counter[0] ;
 wire \u_window_buffer.read_ptr[0] ;
 wire \u_window_buffer.read_ptr[10] ;
 wire \u_window_buffer.read_ptr[11] ;
 wire \u_window_buffer.read_ptr[12] ;
 wire \u_window_buffer.read_ptr[13] ;
 wire \u_window_buffer.read_ptr[14] ;
 wire \u_window_buffer.read_ptr[15] ;
 wire \u_window_buffer.read_ptr[16] ;
 wire \u_window_buffer.read_ptr[17] ;
 wire \u_window_buffer.read_ptr[18] ;
 wire \u_window_buffer.read_ptr[19] ;
 wire \u_window_buffer.read_ptr[1] ;
 wire \u_window_buffer.read_ptr[20] ;
 wire \u_window_buffer.read_ptr[21] ;
 wire \u_window_buffer.read_ptr[22] ;
 wire \u_window_buffer.read_ptr[23] ;
 wire \u_window_buffer.read_ptr[24] ;
 wire \u_window_buffer.read_ptr[25] ;
 wire \u_window_buffer.read_ptr[26] ;
 wire \u_window_buffer.read_ptr[27] ;
 wire \u_window_buffer.read_ptr[28] ;
 wire \u_window_buffer.read_ptr[29] ;
 wire \u_window_buffer.read_ptr[2] ;
 wire \u_window_buffer.read_ptr[30] ;
 wire \u_window_buffer.read_ptr[3] ;
 wire \u_window_buffer.read_ptr[4] ;
 wire \u_window_buffer.read_ptr[5] ;
 wire \u_window_buffer.read_ptr[6] ;
 wire \u_window_buffer.read_ptr[7] ;
 wire \u_window_buffer.read_ptr[8] ;
 wire \u_window_buffer.read_ptr[9] ;
 wire \u_window_buffer.write_ptr[0] ;
 wire \u_window_buffer.write_ptr[1] ;
 wire net2928;
 wire net2927;
 wire net2926;
 wire net2924;
 wire net2923;
 wire net2921;
 wire net2920;
 wire net2918;
 wire net2919;
 wire net2917;
 wire net2916;
 wire net2915;
 wire net2914;
 wire net2912;
 wire net2911;
 wire net2910;
 wire net2908;
 wire net2907;
 wire net2906;
 wire net2905;
 wire net2904;
 wire net2903;
 wire net2902;
 wire net2901;
 wire net2909;
 wire net2900;
 wire net2898;
 wire net2897;
 wire net2896;
 wire net2895;
 wire net2894;
 wire net2893;
 wire net2892;
 wire net2888;
 wire net2887;
 wire net2886;
 wire net2885;
 wire net2884;
 wire net2883;
 wire net2882;
 wire net2880;
 wire net2878;
 wire net2877;
 wire net2874;
 wire net2873;
 wire net2872;
 wire net2871;
 wire net2869;
 wire net2870;
 wire net2867;
 wire net2865;
 wire net2864;
 wire net2866;
 wire net2863;
 wire net2862;
 wire net2861;
 wire net2860;
 wire net2859;
 wire net2868;
 wire net2858;
 wire net2857;
 wire net2854;
 wire net2853;
 wire net2852;
 wire net2855;
 wire net2851;
 wire net2856;
 wire net2850;
 wire net2849;
 wire net2848;
 wire net2847;
 wire net2846;
 wire net2875;
 wire net2843;
 wire net2842;
 wire net2841;
 wire net2840;
 wire net2838;
 wire net2836;
 wire net2835;
 wire net2833;
 wire net2832;
 wire net2831;
 wire net2834;
 wire net2829;
 wire net2828;
 wire net2827;
 wire net2825;
 wire net2824;
 wire net2822;
 wire net2823;
 wire net2821;
 wire net2820;
 wire net2819;
 wire net2817;
 wire net2816;
 wire net2815;
 wire net2814;
 wire net2813;
 wire net2811;
 wire net2810;
 wire net2809;
 wire net2808;
 wire net2807;
 wire net2806;
 wire net2805;
 wire net2804;
 wire net2803;
 wire net2802;
 wire net2800;
 wire net2799;
 wire net2798;
 wire net2797;
 wire net2796;
 wire net2795;
 wire net2794;
 wire net2793;
 wire net2790;
 wire net2789;
 wire net2788;
 wire net2786;
 wire net2785;
 wire net2784;
 wire net2783;
 wire net2782;
 wire net2779;
 wire net2778;
 wire net2777;
 wire net2776;
 wire net2774;
 wire net2773;
 wire net2772;
 wire net2771;
 wire net2769;
 wire net2768;
 wire net2770;
 wire net2767;
 wire net2765;
 wire net2762;
 wire net2760;
 wire net2758;
 wire net2756;
 wire net2755;
 wire net2754;
 wire net2752;
 wire net2751;
 wire net2750;
 wire net2747;
 wire net6028;
 wire net2745;
 wire net2743;
 wire net2742;
 wire net2741;
 wire net5731;
 wire net2740;
 wire net2739;
 wire net2748;
 wire net2738;
 wire net2736;
 wire net2737;
 wire net2733;
 wire net2732;
 wire net2731;
 wire net2730;
 wire net2729;
 wire net5725;
 wire net2727;
 wire net5730;
 wire net2735;
 wire net2734;
 wire net2725;
 wire net2723;
 wire net2722;
 wire net2720;
 wire net2719;
 wire net2718;
 wire net2724;
 wire net2721;
 wire net2715;
 wire net2714;
 wire net6027;
 wire net2711;
 wire net2712;
 wire net2709;
 wire net2708;
 wire net2707;
 wire net2706;
 wire net2704;
 wire net2713;
 wire net2710;
 wire net2703;
 wire net2705;
 wire net2699;
 wire net2697;
 wire net2700;
 wire net2698;
 wire net2696;
 wire net2702;
 wire clknet_leaf_1_clk;
 wire net2701;
 wire clknet_leaf_0_clk;
 wire net2717;
 wire net2716;
 wire net212;
 wire net211;
 wire net210;
 wire net209;
 wire net3056;
 wire net3057;
 wire net3061;
 wire net3060;
 wire net3062;
 wire net3089;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3156;
 wire net3155;
 wire net3132;
 wire net3133;
 wire net3142;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3147;
 wire net3146;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3150;
 wire net3148;
 wire net3149;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3190;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3198;
 wire net3199;
 wire net3211;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3208;
 wire net3207;
 wire net3209;
 wire net3210;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3225;
 wire net3223;
 wire net3224;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3230;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3243;
 wire net3245;
 wire net3255;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3256;
 wire net3257;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3266;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3281;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3294;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3322;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3318;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3323;
 wire net3324;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3332;
 wire net3334;
 wire net3343;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3344;
 wire net3453;
 wire net3345;
 wire net3349;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3448;
 wire net3378;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3430;
 wire net3379;
 wire net3380;
 wire net3425;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3400;
 wire net3399;
 wire net3422;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3408;
 wire net3406;
 wire net3407;
 wire net3418;
 wire net3409;
 wire net3413;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3423;
 wire net3424;
 wire net3426;
 wire net3427;
 wire net5910;
 wire net3429;
 wire net3440;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3533;
 wire net3513;
 wire net3506;
 wire net3463;
 wire net3482;
 wire net3469;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3497;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3512;
 wire net3511;
 wire net3518;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3534;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3560;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net6001;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3591;
 wire net3592;
 wire net3613;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3603;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3609;
 wire net3607;
 wire net3608;
 wire net3611;
 wire net3610;
 wire net3612;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3634;
 wire net3639;
 wire net3637;
 wire net3638;
 wire net3640;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3647;
 wire net6002;
 wire net3649;
 wire net3656;
 wire net3650;
 wire net3651;
 wire net3652;
 wire net3655;
 wire net3653;
 wire net3654;
 wire net3657;
 wire net3658;
 wire net3670;
 wire net3660;
 wire net3661;
 wire net3662;
 wire net3668;
 wire net3663;
 wire net3664;
 wire net3665;
 wire net3666;
 wire net3667;
 wire net3669;
 wire net3671;
 wire net3672;
 wire net3673;
 wire net3674;
 wire net3675;
 wire net3676;
 wire net3681;
 wire net3678;
 wire net3679;
 wire net3680;
 wire net3682;
 wire net3683;
 wire net3684;
 wire net3703;
 wire net3685;
 wire net3686;
 wire net3687;
 wire net3702;
 wire net3688;
 wire net3694;
 wire net3689;
 wire net3690;
 wire net3691;
 wire net3692;
 wire net3693;
 wire net3695;
 wire net3696;
 wire net3697;
 wire net3698;
 wire net3699;
 wire net3700;
 wire net3701;
 wire net3704;
 wire net3706;
 wire net3708;
 wire net3709;
 wire net3710;
 wire net3712;
 wire net3716;
 wire net3717;
 wire net3718;
 wire net3723;
 wire net3719;
 wire net3720;
 wire net3721;
 wire net3722;
 wire net3724;
 wire net3726;
 wire net3729;
 wire net3728;
 wire net3731;
 wire net3730;
 wire net3732;
 wire net3733;
 wire net3735;
 wire net3736;
 wire net3737;
 wire net3738;
 wire net3739;
 wire net3740;
 wire net3741;
 wire net3742;
 wire net3743;
 wire net3744;
 wire net3745;
 wire net3746;
 wire net3747;
 wire net3753;
 wire net3748;
 wire net3749;
 wire net3750;
 wire net3751;
 wire net3752;
 wire net3766;
 wire net3764;
 wire net3756;
 wire net3757;
 wire net3758;
 wire net3759;
 wire net3760;
 wire net3761;
 wire net3762;
 wire net3763;
 wire net3765;
 wire net3767;
 wire net3768;
 wire net3769;
 wire net3774;
 wire net3771;
 wire net3772;
 wire net3773;
 wire net3775;
 wire net3782;
 wire net3778;
 wire net3777;
 wire net3779;
 wire net3780;
 wire net3781;
 wire net3783;
 wire net3784;
 wire net3785;
 wire net3786;
 wire net3787;
 wire net3789;
 wire net3791;
 wire net3792;
 wire net3798;
 wire net3794;
 wire net3795;
 wire net3796;
 wire net3797;
 wire net3799;
 wire net3800;
 wire net3801;
 wire net3802;
 wire net3803;
 wire net3804;
 wire net3805;
 wire net3806;
 wire net3807;
 wire net3809;
 wire net3811;
 wire net3813;
 wire net3814;
 wire net3815;
 wire net3816;
 wire net3817;
 wire net3818;
 wire net3819;
 wire net3820;
 wire net3824;
 wire net3823;
 wire net3825;
 wire net3827;
 wire net3828;
 wire net3829;
 wire net3878;
 wire net3830;
 wire net3831;
 wire net3832;
 wire net3833;
 wire net3841;
 wire net3834;
 wire net3835;
 wire net3836;
 wire net3837;
 wire net3838;
 wire net3839;
 wire net3840;
 wire net3848;
 wire net3842;
 wire net3843;
 wire net3844;
 wire net3845;
 wire net3846;
 wire net3847;
 wire net3858;
 wire net3849;
 wire net3850;
 wire net3851;
 wire net3852;
 wire net3853;
 wire net3854;
 wire net3855;
 wire net3856;
 wire net3857;
 wire net3859;
 wire net3860;
 wire net3861;
 wire net3862;
 wire net3863;
 wire net3869;
 wire net3864;
 wire net3865;
 wire net3866;
 wire net3867;
 wire net3868;
 wire net3870;
 wire net3871;
 wire net3872;
 wire net3873;
 wire net3874;
 wire net3875;
 wire net3876;
 wire net3877;
 wire net3881;
 wire net3879;
 wire net3880;
 wire net3913;
 wire net3882;
 wire net3883;
 wire net3884;
 wire net3889;
 wire net3885;
 wire net3886;
 wire net3887;
 wire net3888;
 wire net3890;
 wire net3891;
 wire net3892;
 wire net3893;
 wire net3894;
 wire net3895;
 wire net3896;
 wire net3897;
 wire net3901;
 wire net3898;
 wire net3899;
 wire net3900;
 wire net3902;
 wire net3903;
 wire net3904;
 wire net3905;
 wire net3906;
 wire net3907;
 wire net3908;
 wire net3909;
 wire net3910;
 wire net3912;
 wire net3911;
 wire net3914;
 wire net3915;
 wire net3916;
 wire net3920;
 wire net3917;
 wire net3918;
 wire net3919;
 wire net3921;
 wire net3923;
 wire net3924;
 wire net3925;
 wire net3926;
 wire net3928;
 wire net3929;
 wire net3930;
 wire net3932;
 wire net3933;
 wire net3935;
 wire net3939;
 wire net3936;
 wire net3937;
 wire net3938;
 wire net3941;
 wire net3942;
 wire net3943;
 wire net3944;
 wire net3945;
 wire net3946;
 wire net3947;
 wire net3948;
 wire net3949;
 wire net3950;
 wire net3951;
 wire net3952;
 wire net3954;
 wire net3955;
 wire net3956;
 wire net3979;
 wire net3957;
 wire net3958;
 wire net3959;
 wire net3960;
 wire net3965;
 wire net3961;
 wire net3962;
 wire net3963;
 wire net3964;
 wire net3974;
 wire net3966;
 wire net3967;
 wire net3968;
 wire net3969;
 wire net3973;
 wire net3970;
 wire net3971;
 wire net3972;
 wire net3975;
 wire net3976;
 wire net3977;
 wire net3978;
 wire net3980;
 wire net3981;
 wire net3982;
 wire net3985;
 wire net3986;
 wire net3987;
 wire net3989;
 wire net3990;
 wire net3991;
 wire net4028;
 wire net3992;
 wire net4021;
 wire net3993;
 wire net3994;
 wire net3999;
 wire net3995;
 wire net3996;
 wire net3997;
 wire net3998;
 wire net4020;
 wire net4000;
 wire net4018;
 wire net4016;
 wire net4008;
 wire net4004;
 wire net4017;
 wire net4001;
 wire net4002;
 wire net4003;
 wire net4005;
 wire net4006;
 wire net4007;
 wire net4010;
 wire net4009;
 wire net4011;
 wire net4012;
 wire net4013;
 wire net4014;
 wire net4015;
 wire net4019;
 wire net4022;
 wire net4023;
 wire net4024;
 wire net4025;
 wire net4026;
 wire net4027;
 wire net4029;
 wire net4030;
 wire net4031;
 wire net4032;
 wire net4037;
 wire net4033;
 wire net4034;
 wire net4035;
 wire net4036;
 wire net4038;
 wire net4039;
 wire net4040;
 wire net4043;
 wire net4042;
 wire net4044;
 wire net4045;
 wire net4046;
 wire net4047;
 wire net4048;
 wire net4049;
 wire net4050;
 wire net4051;
 wire net4064;
 wire net4053;
 wire net4054;
 wire net4055;
 wire net4056;
 wire net4057;
 wire net4061;
 wire net4058;
 wire net4059;
 wire net4060;
 wire net4062;
 wire net4063;
 wire net4066;
 wire net4067;
 wire net4068;
 wire net4070;
 wire net4071;
 wire net4072;
 wire net4073;
 wire net4074;
 wire net4084;
 wire net4076;
 wire net4077;
 wire net4078;
 wire net4079;
 wire net4080;
 wire net4081;
 wire net4082;
 wire net4083;
 wire net4085;
 wire net4087;
 wire net4088;
 wire net4089;
 wire net4090;
 wire net4091;
 wire net4092;
 wire net4093;
 wire net4094;
 wire net4095;
 wire net4096;
 wire net4097;
 wire net4098;
 wire net4099;
 wire net4100;
 wire net4101;
 wire net4102;
 wire net4103;
 wire net4104;
 wire net4105;
 wire net4108;
 wire net4110;
 wire net4109;
 wire net4114;
 wire net4111;
 wire net4112;
 wire net4113;
 wire net4122;
 wire net4115;
 wire net4116;
 wire net4117;
 wire net4118;
 wire net4119;
 wire net4120;
 wire net4121;
 wire net4123;
 wire net4124;
 wire net4126;
 wire net4127;
 wire net4130;
 wire net4129;
 wire net4131;
 wire net4132;
 wire net4134;
 wire net4136;
 wire net4135;
 wire net4143;
 wire net4137;
 wire net4138;
 wire net4139;
 wire net4140;
 wire net4141;
 wire net4142;
 wire net4144;
 wire net4145;
 wire net4146;
 wire net4148;
 wire net4149;
 wire net4150;
 wire net4151;
 wire net4152;
 wire net4153;
 wire net4154;
 wire net4155;
 wire net4156;
 wire net4158;
 wire net4159;
 wire net4161;
 wire net4164;
 wire net4165;
 wire net4166;
 wire net4168;
 wire net4171;
 wire net4170;
 wire net4172;
 wire net4173;
 wire net4174;
 wire net4175;
 wire net4176;
 wire net4177;
 wire net4178;
 wire net4179;
 wire net4180;
 wire net4189;
 wire net4182;
 wire net4183;
 wire net4184;
 wire net4185;
 wire net4186;
 wire net4187;
 wire net4188;
 wire net4190;
 wire net4191;
 wire net4192;
 wire net4193;
 wire net4194;
 wire net4196;
 wire net4195;
 wire net4210;
 wire net4197;
 wire net4198;
 wire net4199;
 wire net4200;
 wire net4201;
 wire net4207;
 wire net4203;
 wire net4202;
 wire net4204;
 wire net4205;
 wire net4206;
 wire net4208;
 wire net4209;
 wire net4211;
 wire net4212;
 wire net4246;
 wire net4213;
 wire net4214;
 wire net4236;
 wire net4215;
 wire net4216;
 wire net4217;
 wire net4228;
 wire net4218;
 wire net4219;
 wire net4220;
 wire net4221;
 wire net4222;
 wire net4223;
 wire net4224;
 wire net4225;
 wire net4226;
 wire net4227;
 wire net4229;
 wire net4230;
 wire net4231;
 wire net4232;
 wire net4233;
 wire net4234;
 wire net4235;
 wire net4237;
 wire net4238;
 wire net4239;
 wire net4240;
 wire net4242;
 wire net4241;
 wire net4243;
 wire net4244;
 wire net4245;
 wire net4255;
 wire net4247;
 wire net4248;
 wire net4249;
 wire net4250;
 wire net4251;
 wire net4252;
 wire net4253;
 wire net4254;
 wire net4257;
 wire net4256;
 wire net4262;
 wire net4263;
 wire net4264;
 wire net4265;
 wire net4266;
 wire net4276;
 wire net4267;
 wire net4268;
 wire net4269;
 wire net4270;
 wire net4271;
 wire net4272;
 wire net4273;
 wire net4274;
 wire net4275;
 wire net4287;
 wire net4277;
 wire net4285;
 wire net4278;
 wire net4279;
 wire net4280;
 wire net4281;
 wire net4282;
 wire net4283;
 wire net4284;
 wire net4286;
 wire net4307;
 wire net4297;
 wire net4294;
 wire net4292;
 wire net4291;
 wire net4293;
 wire net4295;
 wire net4296;
 wire net4301;
 wire net4298;
 wire net4299;
 wire net4300;
 wire net4306;
 wire net4303;
 wire net4302;
 wire net4304;
 wire net4305;
 wire net4308;
 wire net4309;
 wire net4311;
 wire net4312;
 wire net4313;
 wire net4314;
 wire net4315;
 wire net4316;
 wire net4317;
 wire net4318;
 wire net4341;
 wire net4330;
 wire net4319;
 wire net4320;
 wire net4321;
 wire net4322;
 wire net4329;
 wire net4323;
 wire net4324;
 wire net4325;
 wire net4326;
 wire net4327;
 wire net4328;
 wire net4331;
 wire net4332;
 wire net4333;
 wire net4334;
 wire net4335;
 wire net4336;
 wire net4337;
 wire net4338;
 wire net4339;
 wire net4340;
 wire net4343;
 wire net4344;
 wire net4348;
 wire net4345;
 wire net4346;
 wire net4347;
 wire net4350;
 wire net4351;
 wire net4352;
 wire net4354;
 wire net4362;
 wire net4356;
 wire net4357;
 wire net4358;
 wire net4359;
 wire net4360;
 wire net4361;
 wire net4369;
 wire net4364;
 wire net4365;
 wire net4366;
 wire net4367;
 wire net4368;
 wire net4370;
 wire net4371;
 wire net4372;
 wire net4373;
 wire net4374;
 wire net4375;
 wire net4376;
 wire net4377;
 wire net4378;
 wire net4379;
 wire net4380;
 wire net4381;
 wire net4392;
 wire net4382;
 wire net4383;
 wire net4384;
 wire net4385;
 wire net4386;
 wire net4387;
 wire net4389;
 wire net4388;
 wire net4390;
 wire net4391;
 wire net4393;
 wire net4394;
 wire net4395;
 wire net4396;
 wire net4398;
 wire net4399;
 wire net4400;
 wire net4424;
 wire net4409;
 wire net4403;
 wire net4404;
 wire net4405;
 wire net4406;
 wire net4407;
 wire net4408;
 wire net4421;
 wire net4410;
 wire net4411;
 wire net4412;
 wire net4413;
 wire net4414;
 wire net4415;
 wire net4416;
 wire net4417;
 wire net4418;
 wire net4419;
 wire net4420;
 wire net4422;
 wire net4423;
 wire net4426;
 wire net4428;
 wire net4429;
 wire net4446;
 wire net4432;
 wire net4442;
 wire net4433;
 wire net4434;
 wire net4435;
 wire net4436;
 wire net4437;
 wire net4438;
 wire net4439;
 wire net4440;
 wire net4441;
 wire net4443;
 wire net4444;
 wire net4445;
 wire net4592;
 wire net4447;
 wire net4448;
 wire net4460;
 wire net4450;
 wire net4449;
 wire net4451;
 wire net4452;
 wire net4456;
 wire net4453;
 wire net4454;
 wire net4455;
 wire net4457;
 wire net4458;
 wire net4459;
 wire net4586;
 wire net4464;
 wire net4461;
 wire net4462;
 wire net4463;
 wire net4585;
 wire net4465;
 wire net4466;
 wire net4467;
 wire net4468;
 wire net4469;
 wire net4581;
 wire net4470;
 wire net4471;
 wire net4472;
 wire net4575;
 wire net4473;
 wire net4474;
 wire net4475;
 wire net4476;
 wire net4570;
 wire net4477;
 wire net4478;
 wire net4479;
 wire net4560;
 wire net4480;
 wire net4481;
 wire net4528;
 wire net4482;
 wire net4506;
 wire net4483;
 wire net4484;
 wire net4485;
 wire net4486;
 wire net4487;
 wire net4488;
 wire net4489;
 wire net4490;
 wire net4491;
 wire net4492;
 wire net4493;
 wire net4494;
 wire net4502;
 wire net4495;
 wire net4496;
 wire net4497;
 wire net4499;
 wire net4498;
 wire net4500;
 wire net4501;
 wire net4503;
 wire net4504;
 wire net4505;
 wire net4507;
 wire net4508;
 wire net4509;
 wire net4510;
 wire net4511;
 wire net4512;
 wire net4513;
 wire net4514;
 wire net4515;
 wire net4516;
 wire net4517;
 wire net4518;
 wire net4523;
 wire net4519;
 wire net4520;
 wire net4521;
 wire net4522;
 wire net4524;
 wire net4525;
 wire net4526;
 wire net4527;
 wire net4559;
 wire net4529;
 wire net4530;
 wire net4531;
 wire net4532;
 wire net4533;
 wire net4534;
 wire net4535;
 wire net4536;
 wire net4537;
 wire net4538;
 wire net4541;
 wire net4539;
 wire net4540;
 wire net4542;
 wire net4558;
 wire net4543;
 wire net4544;
 wire net4557;
 wire net4545;
 wire net4546;
 wire net4547;
 wire net4548;
 wire net4549;
 wire net4550;
 wire net4551;
 wire net4552;
 wire net4553;
 wire net4554;
 wire net4555;
 wire net4556;
 wire net4561;
 wire net4562;
 wire net4563;
 wire net4564;
 wire net4565;
 wire net4566;
 wire net4567;
 wire net4568;
 wire net4569;
 wire net4573;
 wire net4571;
 wire net4572;
 wire net4574;
 wire net4576;
 wire net4577;
 wire net4580;
 wire net4578;
 wire net4579;
 wire net4582;
 wire net4583;
 wire net4584;
 wire net4587;
 wire net4588;
 wire net4589;
 wire net4590;
 wire net4591;
 wire net4596;
 wire net4655;
 wire net4597;
 wire net4598;
 wire net4599;
 wire net4635;
 wire net4634;
 wire net4633;
 wire net4600;
 wire net4601;
 wire net4602;
 wire net4603;
 wire net4632;
 wire net4604;
 wire net4605;
 wire net4609;
 wire net4606;
 wire net4607;
 wire net4608;
 wire net4610;
 wire net4611;
 wire net4612;
 wire net4631;
 wire net4630;
 wire net4613;
 wire net4614;
 wire net4615;
 wire net4616;
 wire net4617;
 wire net4618;
 wire net4619;
 wire net4620;
 wire net4621;
 wire net4622;
 wire net4627;
 wire net4623;
 wire net4626;
 wire net4624;
 wire net4625;
 wire net4628;
 wire net4629;
 wire net4649;
 wire net4641;
 wire net4639;
 wire net4637;
 wire net4636;
 wire net4647;
 wire net4638;
 wire net4640;
 wire net4642;
 wire net4643;
 wire net4646;
 wire net4644;
 wire net4645;
 wire net4648;
 wire net4651;
 wire net4650;
 wire net4653;
 wire net4652;
 wire net4654;
 wire net5033;
 wire net5032;
 wire net5027;
 wire net4657;
 wire net4696;
 wire net4695;
 wire net4694;
 wire net4693;
 wire net4674;
 wire net4662;
 wire net4658;
 wire net4659;
 wire net4660;
 wire net4661;
 wire net4663;
 wire net4664;
 wire net4665;
 wire net4666;
 wire net4667;
 wire net4668;
 wire net4669;
 wire net4670;
 wire net4671;
 wire net4672;
 wire net4673;
 wire net4683;
 wire net4675;
 wire net4676;
 wire net4677;
 wire net4678;
 wire net4679;
 wire net4680;
 wire net4681;
 wire net4682;
 wire net4689;
 wire net4684;
 wire net4685;
 wire net4686;
 wire net4687;
 wire net4688;
 wire net4690;
 wire net4691;
 wire net4692;
 wire net5026;
 wire net4697;
 wire net4698;
 wire net4699;
 wire net4700;
 wire net4701;
 wire net5025;
 wire net5024;
 wire net4708;
 wire net4702;
 wire net4703;
 wire net4704;
 wire net4705;
 wire net4706;
 wire net4707;
 wire net4709;
 wire net4710;
 wire net5023;
 wire net5011;
 wire net5000;
 wire net4998;
 wire net4921;
 wire net4920;
 wire net4915;
 wire net4904;
 wire net4902;
 wire net4901;
 wire net4900;
 wire net4711;
 wire net4712;
 wire net4713;
 wire net4899;
 wire net4716;
 wire net4715;
 wire net4714;
 wire net4898;
 wire net4891;
 wire net4894;
 wire net4890;
 wire net4888;
 wire net4761;
 wire net4758;
 wire net4754;
 wire net4751;
 wire net4749;
 wire net4747;
 wire net4740;
 wire net4739;
 wire net4737;
 wire net4735;
 wire net4727;
 wire net4717;
 wire net4724;
 wire net4719;
 wire net4718;
 wire net4720;
 wire net4721;
 wire net4722;
 wire net4723;
 wire net4725;
 wire net4726;
 wire net4728;
 wire net4729;
 wire net4730;
 wire net4731;
 wire net4732;
 wire net4733;
 wire net4734;
 wire net4736;
 wire net4738;
 wire net4741;
 wire net4742;
 wire net4743;
 wire net4744;
 wire net4745;
 wire net4746;
 wire net4748;
 wire net4750;
 wire net4752;
 wire net4753;
 wire net4755;
 wire net4756;
 wire net4757;
 wire net4760;
 wire net4759;
 wire net4884;
 wire net4762;
 wire net4871;
 wire net4764;
 wire net4763;
 wire net4868;
 wire net4801;
 wire net4765;
 wire net4768;
 wire net4766;
 wire net4767;
 wire net4770;
 wire net4769;
 wire net4772;
 wire net4771;
 wire net4774;
 wire net4773;
 wire net4776;
 wire net4775;
 wire net4778;
 wire net4777;
 wire net4780;
 wire net4779;
 wire net4782;
 wire net4781;
 wire net4784;
 wire net4783;
 wire net4786;
 wire net4785;
 wire net4788;
 wire net4787;
 wire net4790;
 wire net4789;
 wire net4792;
 wire net4791;
 wire net4794;
 wire net4793;
 wire net4796;
 wire net4795;
 wire net4798;
 wire net4797;
 wire net4800;
 wire net4799;
 wire net4803;
 wire net4802;
 wire net4805;
 wire net4804;
 wire net4807;
 wire net4806;
 wire net4865;
 wire net4809;
 wire net4808;
 wire net4811;
 wire net4810;
 wire net4864;
 wire net4860;
 wire net4812;
 wire net4851;
 wire net4813;
 wire net4850;
 wire net4848;
 wire net4814;
 wire net4815;
 wire net4816;
 wire net4817;
 wire net4818;
 wire net4819;
 wire net4820;
 wire net4821;
 wire net4822;
 wire net4823;
 wire net4824;
 wire net4826;
 wire net4825;
 wire net4846;
 wire net4827;
 wire net4828;
 wire net4840;
 wire net4839;
 wire net4829;
 wire net4830;
 wire net4833;
 wire net4831;
 wire net4832;
 wire net4835;
 wire net4834;
 wire net4836;
 wire net4837;
 wire net4838;
 wire net4841;
 wire net4842;
 wire net4844;
 wire net4843;
 wire net4845;
 wire net4847;
 wire net4849;
 wire net4852;
 wire net4853;
 wire net4858;
 wire net4854;
 wire net4855;
 wire net4856;
 wire net4857;
 wire net4859;
 wire net4861;
 wire net4862;
 wire net4863;
 wire net4866;
 wire net4867;
 wire net4869;
 wire net4870;
 wire net4883;
 wire net4872;
 wire net4873;
 wire net4874;
 wire net4875;
 wire net4876;
 wire net4877;
 wire net4878;
 wire net4880;
 wire net4879;
 wire net4881;
 wire net4882;
 wire net4885;
 wire net4886;
 wire net4887;
 wire net4889;
 wire net4892;
 wire net4893;
 wire net4895;
 wire net4896;
 wire net4897;
 wire net4903;
 wire net4905;
 wire net4906;
 wire net4907;
 wire net4908;
 wire net4909;
 wire net4910;
 wire net4911;
 wire net4912;
 wire net4913;
 wire net4914;
 wire net4916;
 wire net4917;
 wire net4918;
 wire net4919;
 wire net4925;
 wire net4922;
 wire net4923;
 wire net4924;
 wire net4926;
 wire net4927;
 wire net4928;
 wire net4929;
 wire net4930;
 wire net4931;
 wire net4997;
 wire net4932;
 wire net4935;
 wire net4933;
 wire net4934;
 wire net4936;
 wire net4937;
 wire net4938;
 wire net4939;
 wire net4940;
 wire net4941;
 wire net4942;
 wire net4943;
 wire net4944;
 wire net4945;
 wire net4946;
 wire net4947;
 wire net4948;
 wire net4949;
 wire net4950;
 wire net4951;
 wire net4952;
 wire net4953;
 wire net4954;
 wire net4955;
 wire net4956;
 wire net4957;
 wire net4958;
 wire net4959;
 wire net4960;
 wire net4961;
 wire net4962;
 wire net4963;
 wire net4964;
 wire net4965;
 wire net4966;
 wire net4967;
 wire net4968;
 wire net4969;
 wire net4970;
 wire net4971;
 wire net4972;
 wire net4973;
 wire net4974;
 wire net4975;
 wire net4976;
 wire net4977;
 wire net4978;
 wire net4979;
 wire net4980;
 wire net4981;
 wire net4982;
 wire net4983;
 wire net4984;
 wire net4985;
 wire net4986;
 wire net4987;
 wire net4988;
 wire net4989;
 wire net4990;
 wire net4991;
 wire net4992;
 wire net4993;
 wire net4994;
 wire net4995;
 wire net4996;
 wire net4999;
 wire net5001;
 wire net5002;
 wire net5003;
 wire net5004;
 wire net5005;
 wire net5006;
 wire net5007;
 wire net5008;
 wire net5009;
 wire net5010;
 wire net5012;
 wire net5013;
 wire net5014;
 wire net5015;
 wire net5016;
 wire net5017;
 wire net5018;
 wire net5019;
 wire net5020;
 wire net5021;
 wire net5022;
 wire net5031;
 wire net5030;
 wire net5029;
 wire net5028;
 wire net5044;
 wire net5040;
 wire net5035;
 wire net5034;
 wire net5036;
 wire net5037;
 wire net5038;
 wire net5039;
 wire net5041;
 wire net5043;
 wire net5042;
 wire net5045;
 wire net5046;
 wire net5047;
 wire net5048;
 wire net5056;
 wire net5057;
 wire net5058;
 wire net5061;
 wire net5064;
 wire net5065;
 wire net5066;
 wire net5067;
 wire net5068;
 wire net5083;
 wire net5070;
 wire net5071;
 wire net5072;
 wire net5073;
 wire net5074;
 wire net5075;
 wire net5076;
 wire net5077;
 wire net5078;
 wire net5082;
 wire net5079;
 wire net5080;
 wire net5081;
 wire net5084;
 wire net5085;
 wire net5086;
 wire net5087;
 wire net5093;
 wire net5089;
 wire net5090;
 wire net5091;
 wire net5092;
 wire net5190;
 wire net5094;
 wire net5098;
 wire net5095;
 wire net5096;
 wire net5097;
 wire net5099;
 wire net5100;
 wire net5111;
 wire net5101;
 wire net5102;
 wire net5103;
 wire net5104;
 wire net5105;
 wire net5106;
 wire net5107;
 wire net5108;
 wire net5109;
 wire net5110;
 wire net5112;
 wire net5113;
 wire net5114;
 wire net5115;
 wire net5116;
 wire net5117;
 wire net5118;
 wire net5119;
 wire net5120;
 wire net5121;
 wire net5122;
 wire net5123;
 wire net5124;
 wire net5125;
 wire net5126;
 wire net5127;
 wire net5128;
 wire net5129;
 wire net5130;
 wire net5131;
 wire net5132;
 wire net5133;
 wire net5134;
 wire net5135;
 wire net5136;
 wire net5137;
 wire net5138;
 wire net5139;
 wire net5140;
 wire net5141;
 wire net5142;
 wire net5143;
 wire net5144;
 wire net5145;
 wire net5146;
 wire net5147;
 wire net5148;
 wire net5149;
 wire net5150;
 wire net5151;
 wire net5173;
 wire net5152;
 wire net5153;
 wire net5154;
 wire net5155;
 wire net5156;
 wire net5157;
 wire net5158;
 wire net5162;
 wire net5159;
 wire net5160;
 wire net5161;
 wire net5163;
 wire net5170;
 wire net5164;
 wire net5165;
 wire net5166;
 wire net5167;
 wire net5168;
 wire net5169;
 wire net5171;
 wire net5172;
 wire net5174;
 wire net5175;
 wire net5176;
 wire net5177;
 wire net5178;
 wire net5179;
 wire net5180;
 wire net5181;
 wire net5182;
 wire net5183;
 wire net5184;
 wire net5185;
 wire net5186;
 wire net5187;
 wire net5188;
 wire net5189;
 wire net5191;
 wire net5192;
 wire net5193;
 wire net5194;
 wire net5195;
 wire net5196;
 wire net5197;
 wire net5198;
 wire net5199;
 wire net5201;
 wire net5202;
 wire net5203;
 wire net5204;
 wire net5205;
 wire net5211;
 wire net5206;
 wire net5207;
 wire net5208;
 wire net5209;
 wire net5210;
 wire net5212;
 wire net5227;
 wire net5213;
 wire net5214;
 wire net5215;
 wire net5216;
 wire net5217;
 wire net5218;
 wire net5219;
 wire net5220;
 wire net5221;
 wire net5222;
 wire net5223;
 wire net5224;
 wire net5225;
 wire net5226;
 wire net5229;
 wire net5230;
 wire net5231;
 wire net5232;
 wire net5233;
 wire net5234;
 wire net5237;
 wire net5238;
 wire net5239;
 wire net5240;
 wire net5253;
 wire net5241;
 wire net5242;
 wire net5251;
 wire net5243;
 wire net5244;
 wire net5245;
 wire net5246;
 wire net5247;
 wire net5248;
 wire net5249;
 wire net5250;
 wire net5252;
 wire net5255;
 wire net5256;
 wire net5257;
 wire net5258;
 wire net5259;
 wire net5261;
 wire net5262;
 wire net5263;
 wire net5264;
 wire net5265;
 wire net5266;
 wire net5267;
 wire net5268;
 wire net5269;
 wire net5270;
 wire net5271;
 wire net5272;
 wire net5273;
 wire net5274;
 wire net5275;
 wire net5276;
 wire net5277;
 wire net5282;
 wire net5278;
 wire net5279;
 wire net5280;
 wire net5281;
 wire net5284;
 wire net5285;
 wire net5286;
 wire net5288;
 wire net5290;
 wire net5293;
 wire net5294;
 wire net5295;
 wire net5296;
 wire net5297;
 wire net5299;
 wire net5298;
 wire net5301;
 wire net5302;
 wire net5303;
 wire net5304;
 wire net5305;
 wire net5306;
 wire net5307;
 wire net5308;
 wire net5309;
 wire net5310;
 wire net5311;
 wire net5312;
 wire net5313;
 wire net5314;
 wire net5315;
 wire net5316;
 wire net5317;
 wire net5318;
 wire net5319;
 wire net5320;
 wire net5321;
 wire net5322;
 wire net5323;
 wire net5324;
 wire net5325;
 wire net5326;
 wire net5328;
 wire net5329;
 wire net5331;
 wire net5332;
 wire net5360;
 wire net5333;
 wire net5334;
 wire net5335;
 wire net5346;
 wire net5336;
 wire net5337;
 wire net5338;
 wire net5339;
 wire net5340;
 wire net5341;
 wire net5342;
 wire net5343;
 wire net5344;
 wire net5345;
 wire net5347;
 wire net5359;
 wire net5348;
 wire net5349;
 wire net5350;
 wire net5351;
 wire net5352;
 wire net5353;
 wire net5354;
 wire net5355;
 wire net5356;
 wire net5357;
 wire net5358;
 wire clknet_leaf_2_clk;
 wire net5363;
 wire net5362;
 wire net2753;
 wire net2757;
 wire net2759;
 wire net2761;
 wire net2763;
 wire net2764;
 wire net2766;
 wire net2775;
 wire net2780;
 wire net2781;
 wire net2787;
 wire net2791;
 wire net2792;
 wire net2801;
 wire net2812;
 wire net2818;
 wire net2826;
 wire net2830;
 wire net2837;
 wire net2839;
 wire net2844;
 wire net2845;
 wire net2876;
 wire net2879;
 wire net2881;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2899;
 wire net2913;
 wire net2922;
 wire net2925;
 wire net2935;
 wire net2943;
 wire net2945;
 wire net2947;
 wire net2948;
 wire net2958;
 wire net2963;
 wire net2967;
 wire net3013;
 wire net3014;
 wire net3059;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3095;
 wire net3101;
 wire net3118;
 wire net3126;
 wire net3130;
 wire net3131;
 wire net3160;
 wire net3161;
 wire net3167;
 wire net3177;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3212;
 wire net3229;
 wire net3231;
 wire net3238;
 wire net3242;
 wire net3244;
 wire net3246;
 wire net3247;
 wire net3258;
 wire net3265;
 wire net3267;
 wire net3276;
 wire net3325;
 wire net3331;
 wire net3333;
 wire net3335;
 wire net3459;
 wire net3535;
 wire net3548;
 wire net3572;
 wire net3576;
 wire net3590;
 wire net3593;
 wire net3618;
 wire net3623;
 wire net3633;
 wire net3635;
 wire net3636;
 wire net3641;
 wire net3646;
 wire net3659;
 wire net3677;
 wire net3705;
 wire net3707;
 wire net3711;
 wire net3713;
 wire net3714;
 wire net3715;
 wire net3725;
 wire net3727;
 wire net3734;
 wire net3754;
 wire net3755;
 wire net3770;
 wire net3776;
 wire net3788;
 wire net3790;
 wire net3793;
 wire net3808;
 wire net3810;
 wire net3812;
 wire net3821;
 wire net3822;
 wire net3826;
 wire net3922;
 wire net3927;
 wire net3931;
 wire net3934;
 wire net3940;
 wire net3953;
 wire net3983;
 wire net3984;
 wire net3988;
 wire net4041;
 wire net4052;
 wire net4065;
 wire net4069;
 wire net4075;
 wire net4086;
 wire net4106;
 wire net4107;
 wire net4125;
 wire net4128;
 wire net4133;
 wire net4147;
 wire net4157;
 wire net4160;
 wire net4162;
 wire net4163;
 wire net4167;
 wire net4169;
 wire net4181;
 wire net4258;
 wire net4259;
 wire net4260;
 wire net4261;
 wire net4288;
 wire net4289;
 wire net4290;
 wire net4310;
 wire net4342;
 wire net4349;
 wire net4353;
 wire net4355;
 wire net4363;
 wire net4397;
 wire net4401;
 wire net4402;
 wire net4425;
 wire net4427;
 wire net4430;
 wire net4431;
 wire net4593;
 wire net4594;
 wire net4595;
 wire net4656;
 wire net5049;
 wire net5050;
 wire net5051;
 wire net5052;
 wire net5053;
 wire net5054;
 wire net5055;
 wire net5059;
 wire net5060;
 wire net5062;
 wire net5063;
 wire net5069;
 wire net5088;
 wire net5200;
 wire net5228;
 wire net5235;
 wire net5236;
 wire net5254;
 wire net5260;
 wire net5283;
 wire net5287;
 wire net5289;
 wire net5291;
 wire net5292;
 wire net5300;
 wire net5327;
 wire net5330;
 wire net5361;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net5364;
 wire net5365;
 wire net5366;
 wire net5367;
 wire net5368;
 wire net5369;
 wire net5370;
 wire net5371;
 wire net5372;
 wire net5373;
 wire net5374;
 wire net5375;
 wire net5376;
 wire net5377;
 wire net5378;
 wire net5379;
 wire net5380;
 wire net5381;
 wire net5382;
 wire net5383;
 wire net5384;
 wire net5385;
 wire net5386;
 wire net5387;
 wire net5388;
 wire net5389;
 wire net5390;
 wire net5391;
 wire net5392;
 wire net5393;
 wire net5394;
 wire net5395;
 wire net5396;
 wire net5397;
 wire net5398;
 wire net5399;
 wire net5400;
 wire net5401;
 wire net5402;
 wire net5403;
 wire net5404;
 wire net5418;
 wire net5419;
 wire net5420;
 wire net5421;
 wire net5422;
 wire net5423;
 wire net5424;
 wire net5425;
 wire net5426;
 wire net5427;
 wire net5428;
 wire net5429;
 wire net5430;
 wire net5431;
 wire net5432;
 wire net5433;
 wire net5434;
 wire net5435;
 wire net5436;
 wire net5437;
 wire net5438;
 wire net5439;
 wire net5440;
 wire net5441;
 wire net5442;
 wire net5443;
 wire net5444;
 wire net5445;
 wire net5446;
 wire net5447;
 wire net5448;
 wire net5449;
 wire net5450;
 wire net5451;
 wire net5452;
 wire net5453;
 wire net5454;
 wire net5455;
 wire net5456;
 wire net5457;
 wire net5458;
 wire net5504;
 wire net5505;
 wire net5506;
 wire net5536;
 wire net5537;
 wire net5538;
 wire net5539;
 wire net5540;
 wire net5541;
 wire net5585;
 wire net5590;
 wire net5591;
 wire net5592;
 wire net5593;
 wire net5594;
 wire net5595;
 wire net5596;
 wire net5597;
 wire net5598;
 wire net5599;
 wire net5600;
 wire net5601;
 wire net5602;
 wire net5603;
 wire net5604;
 wire net5605;
 wire net5606;
 wire net5607;
 wire net5608;
 wire net5609;
 wire net5610;
 wire net5611;
 wire net5612;
 wire net5613;
 wire net5614;
 wire net5615;
 wire net5616;
 wire net5617;
 wire net5618;
 wire net5619;
 wire net5620;
 wire net5621;
 wire net5622;
 wire net5623;
 wire net5624;
 wire net5625;
 wire net5626;
 wire net5627;
 wire net5628;
 wire net5629;
 wire net5630;
 wire net5631;
 wire net5632;
 wire net5633;
 wire net5634;
 wire net5635;
 wire net5636;
 wire net5637;
 wire net5638;
 wire net5653;
 wire net5654;
 wire net5655;
 wire net5661;
 wire net5662;
 wire net5663;
 wire net5664;
 wire net5665;
 wire net5666;
 wire net5667;
 wire net5668;
 wire net5669;
 wire net5670;
 wire net5671;
 wire net5672;
 wire net5673;
 wire net5674;
 wire net5675;
 wire net5676;
 wire net5677;
 wire net5678;
 wire net5679;
 wire net5680;
 wire net5681;
 wire net5682;
 wire net5683;
 wire net5684;
 wire net5685;
 wire net5686;
 wire net5687;
 wire net5688;
 wire net5689;
 wire net5690;
 wire net5691;
 wire net5692;
 wire net5693;
 wire net5694;
 wire net5695;
 wire net5696;
 wire net5697;
 wire net5698;
 wire net5699;
 wire net5700;
 wire net5701;
 wire net5702;
 wire net5703;
 wire net5704;
 wire net5705;
 wire net5706;
 wire net5707;
 wire net5708;
 wire net5709;
 wire net5710;
 wire net5714;
 wire net5715;
 wire net5716;
 wire net5718;
 wire net5719;
 wire net5720;
 wire net5728;
 wire net5757;
 wire net5758;
 wire net5759;
 wire net5760;
 wire net5761;
 wire net5762;
 wire net5763;
 wire net5764;
 wire net5765;
 wire net5766;
 wire net5767;
 wire net5768;
 wire net5769;
 wire net5770;
 wire net5771;
 wire net5772;
 wire net5773;
 wire net5787;
 wire net5819;
 wire net5820;
 wire net5821;
 wire net5822;
 wire net5876;
 wire net5877;
 wire net5887;
 wire net5888;
 wire net5889;
 wire net5894;
 wire net5895;
 wire net5902;
 wire net5903;
 wire net5912;
 wire net5913;
 wire net5914;
 wire net5917;
 wire net5918;
 wire net5920;
 wire net5923;
 wire net5924;
 wire net5933;
 wire net5934;
 wire net5935;
 wire net5936;
 wire net5937;
 wire net5938;
 wire net5939;
 wire net5940;
 wire net5941;
 wire net5957;
 wire net5958;
 wire net5959;
 wire net5960;
 wire net5961;
 wire net5964;
 wire net5972;
 wire net5973;
 wire net5974;
 wire net5975;
 wire net5976;
 wire net5977;
 wire net5978;
 wire net5979;
 wire net5980;
 wire net5981;
 wire net5982;
 wire net5983;
 wire net5984;
 wire net5985;
 wire net5986;
 wire net5987;
 wire net5988;
 wire net5996;
 wire net5997;
 wire net5998;
 wire net5999;
 wire net6000;
 wire net6003;
 wire net6010;
 wire net6011;
 wire net6030;
 wire net6033;
 wire net6034;
 wire net6035;
 wire net6036;
 wire net6037;
 wire net6038;
 wire net6039;
 wire net6040;
 wire net6041;
 wire net6042;
 wire net6043;

 INVx3_ASAP7_75t_R _06546_ (.A(net5363),
    .Y(_06525_));
 BUFx3_ASAP7_75t_R place3055 (.A(_06277_),
    .Y(net3055));
 BUFx3_ASAP7_75t_R place3054 (.A(_02189_),
    .Y(net3054));
 AND3x1_ASAP7_75t_R _06549_ (.A(_00243_),
    .B(_00366_),
    .C(_00365_),
    .Y(_06527_));
 AND3x2_ASAP7_75t_R _06550_ (.A(_06527_),
    .B(_00241_),
    .C(net5279),
    .Y(_06528_));
 AND3x1_ASAP7_75t_R _06551_ (.A(_00237_),
    .B(_00238_),
    .C(_00239_),
    .Y(_00873_));
 AND3x1_ASAP7_75t_R _06552_ (.A(net4866),
    .B(net5277),
    .C(_00873_),
    .Y(_00874_));
 XOR2x2_ASAP7_75t_R _06553_ (.A(_00874_),
    .B(_00236_),
    .Y(_00341_));
 INVx1_ASAP7_75t_R _06554_ (.A(_00242_),
    .Y(_00875_));
 INVx1_ASAP7_75t_R _06555_ (.A(_00243_),
    .Y(_00876_));
 OR3x1_ASAP7_75t_R _06556_ (.A(_00367_),
    .B(_00876_),
    .C(_00875_),
    .Y(_00877_));
 INVx1_ASAP7_75t_R _06557_ (.A(_00877_),
    .Y(_00878_));
 AND3x4_ASAP7_75t_R _06558_ (.A(_00878_),
    .B(_00240_),
    .C(net5278),
    .Y(_00879_));
 AND3x1_ASAP7_75t_R _06559_ (.A(_00879_),
    .B(net5275),
    .C(net5276),
    .Y(_00880_));
 XOR2x2_ASAP7_75t_R _06560_ (.A(_00880_),
    .B(net5274),
    .Y(_00344_));
 AND3x1_ASAP7_75t_R _06561_ (.A(net4866),
    .B(net5276),
    .C(net5277),
    .Y(_00881_));
 XOR2x2_ASAP7_75t_R _06562_ (.A(_00881_),
    .B(net5275),
    .Y(_00347_));
 XOR2x2_ASAP7_75t_R _06563_ (.A(_00879_),
    .B(net5276),
    .Y(_00350_));
 XOR2x2_ASAP7_75t_R _06564_ (.A(_00240_),
    .B(_06528_),
    .Y(_00353_));
 INVx1_ASAP7_75t_R _06565_ (.A(net5278),
    .Y(_00882_));
 XOR2x2_ASAP7_75t_R _06566_ (.A(net4865),
    .B(_00882_),
    .Y(_00356_));
 XOR2x2_ASAP7_75t_R _06567_ (.A(net5082),
    .B(net5279),
    .Y(_00359_));
 XNOR2x2_ASAP7_75t_R _06568_ (.A(net5280),
    .B(net4870),
    .Y(_00362_));
 INVx1_ASAP7_75t_R _06569_ (.A(net5258),
    .Y(\u_fft.sched[45] ));
 INVx1_ASAP7_75t_R _06570_ (.A(_00229_),
    .Y(\u_fft.sched[38] ));
 INVx1_ASAP7_75t_R _06571_ (.A(_00230_),
    .Y(\u_fft.sched[37] ));
 INVx1_ASAP7_75t_R _06572_ (.A(_00231_),
    .Y(\u_fft.sched[36] ));
 INVx1_ASAP7_75t_R _06573_ (.A(_00232_),
    .Y(\u_fft.sched[35] ));
 INVx1_ASAP7_75t_R _06574_ (.A(_00233_),
    .Y(\u_fft.sched[34] ));
 INVx1_ASAP7_75t_R _06575_ (.A(_00234_),
    .Y(\u_fft.sched[33] ));
 INVx1_ASAP7_75t_R _06576_ (.A(_00235_),
    .Y(\u_fft.sched[32] ));
 INVx2_ASAP7_75t_R _06577_ (.A(_00397_),
    .Y(\u_fft.sched[31] ));
 INVx2_ASAP7_75t_R _06578_ (.A(_00396_),
    .Y(\u_fft.sched[30] ));
 OR3x1_ASAP7_75t_R _06579_ (.A(\u_fft.sched[32] ),
    .B(\u_fft.sched[30] ),
    .C(\u_fft.sched[31] ),
    .Y(_00883_));
 OR3x1_ASAP7_75t_R _06580_ (.A(_00883_),
    .B(\u_fft.sched[34] ),
    .C(\u_fft.sched[33] ),
    .Y(_00884_));
 OR3x1_ASAP7_75t_R _06581_ (.A(\u_fft.sched[35] ),
    .B(\u_fft.sched[36] ),
    .C(_00884_),
    .Y(_00885_));
 OR3x1_ASAP7_75t_R _06582_ (.A(\u_fft.sched[37] ),
    .B(\u_fft.sched[38] ),
    .C(_00885_),
    .Y(_00886_));
 XNOR2x2_ASAP7_75t_R _06583_ (.A(_00228_),
    .B(_00886_),
    .Y(_00372_));
 INVx1_ASAP7_75t_R _06584_ (.A(_00398_),
    .Y(_00887_));
 AND3x1_ASAP7_75t_R _06585_ (.A(_00887_),
    .B(net5271),
    .C(net5272),
    .Y(_00888_));
 AND3x1_ASAP7_75t_R _06586_ (.A(_00888_),
    .B(net5269),
    .C(net5270),
    .Y(_00889_));
 AND3x1_ASAP7_75t_R _06587_ (.A(_00889_),
    .B(net5267),
    .C(net5268),
    .Y(_00890_));
 XOR2x2_ASAP7_75t_R _06588_ (.A(_00890_),
    .B(net5078),
    .Y(_00375_));
 XOR2x2_ASAP7_75t_R _06589_ (.A(net4700),
    .B(net5267),
    .Y(_00378_));
 XOR2x2_ASAP7_75t_R _06590_ (.A(_00889_),
    .B(net5076),
    .Y(_00381_));
 XOR2x2_ASAP7_75t_R _06591_ (.A(_00884_),
    .B(net5269),
    .Y(_00384_));
 XOR2x2_ASAP7_75t_R _06592_ (.A(_00888_),
    .B(net5074),
    .Y(_00387_));
 XOR2x2_ASAP7_75t_R _06593_ (.A(net4864),
    .B(net5271),
    .Y(_00390_));
 XOR2x2_ASAP7_75t_R _06594_ (.A(_00398_),
    .B(net5272),
    .Y(_00393_));
 BUFx3_ASAP7_75t_R place3053 (.A(_02196_),
    .Y(net3053));
 INVx1_ASAP7_75t_R _06596_ (.A(net5262),
    .Y(\u_fft.sched[42] ));
 INVx1_ASAP7_75t_R _06597_ (.A(net5263),
    .Y(\u_fft.sched[41] ));
 INVx1_ASAP7_75t_R _06598_ (.A(net5264),
    .Y(\u_fft.sched[40] ));
 BUFx3_ASAP7_75t_R place3052 (.A(_02235_),
    .Y(net3052));
 BUFx3_ASAP7_75t_R place3058 (.A(_06238_),
    .Y(net3058));
 INVx1_ASAP7_75t_R _06601_ (.A(_00332_),
    .Y(_00894_));
 INVx2_ASAP7_75t_R _06602_ (.A(_00164_),
    .Y(_00895_));
 INVx1_ASAP7_75t_R _06603_ (.A(_00165_),
    .Y(_00896_));
 INVx1_ASAP7_75t_R _06604_ (.A(_00329_),
    .Y(_00897_));
 OA21x2_ASAP7_75t_R _06605_ (.A1(_00895_),
    .A2(_00896_),
    .B(_00897_),
    .Y(_00898_));
 INVx1_ASAP7_75t_R _06606_ (.A(net4863),
    .Y(_00899_));
 INVx2_ASAP7_75t_R _06607_ (.A(_00166_),
    .Y(_00900_));
 OR5x1_ASAP7_75t_R _06608_ (.A(_00520_),
    .B(_00900_),
    .C(net5208),
    .D(net5206),
    .E(net5064),
    .Y(_00901_));
 AND2x2_ASAP7_75t_R _06609_ (.A(net5362),
    .B(_00901_),
    .Y(_00902_));
 INVx1_ASAP7_75t_R _06610_ (.A(_00171_),
    .Y(_00903_));
 INVx1_ASAP7_75t_R _06611_ (.A(_00168_),
    .Y(_00904_));
 INVx1_ASAP7_75t_R _06612_ (.A(_00169_),
    .Y(_00905_));
 INVx1_ASAP7_75t_R _06613_ (.A(_00170_),
    .Y(_00906_));
 OR4x1_ASAP7_75t_R _06614_ (.A(_00554_),
    .B(_00905_),
    .C(_00906_),
    .D(_00904_),
    .Y(_00907_));
 INVx1_ASAP7_75t_R _06615_ (.A(_00172_),
    .Y(_00908_));
 INVx1_ASAP7_75t_R _06616_ (.A(_00173_),
    .Y(_00909_));
 INVx1_ASAP7_75t_R _06617_ (.A(_00174_),
    .Y(_00910_));
 OR5x1_ASAP7_75t_R _06618_ (.A(_00907_),
    .B(_00903_),
    .C(_00908_),
    .D(_00909_),
    .E(_00910_),
    .Y(_00911_));
 NOR2x1_ASAP7_75t_R _06619_ (.A(net5205),
    .B(net4751),
    .Y(_00912_));
 AO32x1_ASAP7_75t_R _06620_ (.A1(net5362),
    .A2(net5065),
    .A3(_00899_),
    .B1(_00902_),
    .B2(_00912_),
    .Y(_00015_));
 INVx1_ASAP7_75t_R _06621_ (.A(_00330_),
    .Y(_00913_));
 INVx2_ASAP7_75t_R _06622_ (.A(_00902_),
    .Y(_00914_));
 AO221x1_ASAP7_75t_R _06623_ (.A1(_00322_),
    .A2(_00913_),
    .B1(net5065),
    .B2(net4863),
    .C(_00914_),
    .Y(_00014_));
 AND4x1_ASAP7_75t_R _06624_ (.A(_00205_),
    .B(_00206_),
    .C(_00207_),
    .D(net5243),
    .Y(_00915_));
 AND5x1_ASAP7_75t_R _06625_ (.A(_00201_),
    .B(_00915_),
    .C(_00202_),
    .D(_00203_),
    .E(_00204_),
    .Y(_00916_));
 AND4x1_ASAP7_75t_R _06626_ (.A(_00197_),
    .B(_00198_),
    .C(_00199_),
    .D(_00200_),
    .Y(_00917_));
 AND5x1_ASAP7_75t_R _06627_ (.A(_00193_),
    .B(_00917_),
    .C(net5231),
    .D(_00195_),
    .E(_00196_),
    .Y(_00918_));
 AND3x1_ASAP7_75t_R _06628_ (.A(net5244),
    .B(net5246),
    .C(net5248),
    .Y(_00919_));
 INVx1_ASAP7_75t_R _06629_ (.A(_00550_),
    .Y(_00920_));
 AND5x1_ASAP7_75t_R _06630_ (.A(net5245),
    .B(_00919_),
    .C(_00211_),
    .D(net5247),
    .E(_00920_),
    .Y(_00921_));
 INVx1_ASAP7_75t_R _06631_ (.A(_00190_),
    .Y(_00922_));
 AND4x1_ASAP7_75t_R _06632_ (.A(net5057),
    .B(net5227),
    .C(net5228),
    .D(_00192_),
    .Y(_00923_));
 NOR2x1_ASAP7_75t_R _06633_ (.A(_00186_),
    .B(_00187_),
    .Y(_00924_));
 AND3x1_ASAP7_75t_R _06634_ (.A(net5056),
    .B(net5223),
    .C(net5226),
    .Y(_00925_));
 AND5x1_ASAP7_75t_R _06635_ (.A(_00921_),
    .B(_00918_),
    .C(_00916_),
    .D(_00923_),
    .E(_00925_),
    .Y(_00926_));
 INVx2_ASAP7_75t_R _06636_ (.A(_00926_),
    .Y(_00927_));
 BUFx3_ASAP7_75t_R place3051 (.A(_03912_),
    .Y(net3051));
 INVx1_ASAP7_75t_R _06638_ (.A(_00046_),
    .Y(_00929_));
 NOR2x1_ASAP7_75t_R _06639_ (.A(net5116),
    .B(net5213),
    .Y(_00930_));
 AO21x1_ASAP7_75t_R _06640_ (.A1(net4642),
    .A2(_00929_),
    .B(net5048),
    .Y(_00931_));
 BUFx3_ASAP7_75t_R place3050 (.A(_03916_),
    .Y(net3050));
 BUFx3_ASAP7_75t_R place3049 (.A(_03929_),
    .Y(net3049));
 AND2x2_ASAP7_75t_R _06643_ (.A(_00931_),
    .B(net5363),
    .Y(_00013_));
 INVx1_ASAP7_75t_R _06644_ (.A(_00296_),
    .Y(_00934_));
 INVx1_ASAP7_75t_R _06645_ (.A(_00298_),
    .Y(_00935_));
 OR5x1_ASAP7_75t_R _06646_ (.A(_00295_),
    .B(_00477_),
    .C(_00935_),
    .D(_00297_),
    .E(_00934_),
    .Y(_00936_));
 INVx1_ASAP7_75t_R _06647_ (.A(net5341),
    .Y(_00937_));
 NOR2x1p5_ASAP7_75t_R _06648_ (.A(_00167_),
    .B(_00319_),
    .Y(_00938_));
 AO21x1_ASAP7_75t_R _06649_ (.A1(net5047),
    .A2(_00936_),
    .B(net5046),
    .Y(_00939_));
 BUFx3_ASAP7_75t_R place3047 (.A(_05112_),
    .Y(net3047));
 OR3x1_ASAP7_75t_R _06651_ (.A(_00472_),
    .B(_00300_),
    .C(_00299_),
    .Y(_00941_));
 INVx1_ASAP7_75t_R _06652_ (.A(_00320_),
    .Y(_00942_));
 AND3x1_ASAP7_75t_R _06653_ (.A(_00941_),
    .B(net5362),
    .C(net5045),
    .Y(_00943_));
 AO21x1_ASAP7_75t_R _06654_ (.A1(_00939_),
    .A2(net5362),
    .B(_00943_),
    .Y(_00007_));
 INVx1_ASAP7_75t_R _06655_ (.A(_00167_),
    .Y(_00944_));
 NOR2x1p5_ASAP7_75t_R _06656_ (.A(_00319_),
    .B(_00944_),
    .Y(_00945_));
 BUFx3_ASAP7_75t_R place3046 (.A(_05144_),
    .Y(net3046));
 INVx1_ASAP7_75t_R _06658_ (.A(_00301_),
    .Y(_00947_));
 OR3x1_ASAP7_75t_R _06659_ (.A(net4861),
    .B(net5361),
    .C(_00947_),
    .Y(_00006_));
 INVx1_ASAP7_75t_R _06660_ (.A(net5220),
    .Y(\u_hamming_window.frame_ptr[1] ));
 NOR2x1_ASAP7_75t_R _06661_ (.A(_00046_),
    .B(_00927_),
    .Y(_00948_));
 OR3x1_ASAP7_75t_R _06662_ (.A(_00180_),
    .B(_00181_),
    .C(_00182_),
    .Y(_00949_));
 OR3x1_ASAP7_75t_R _06663_ (.A(_00949_),
    .B(_00024_),
    .C(_00183_),
    .Y(_00950_));
 OR3x1_ASAP7_75t_R _06664_ (.A(_00950_),
    .B(_00178_),
    .C(_00179_),
    .Y(_00951_));
 OR3x1_ASAP7_75t_R _06665_ (.A(net4750),
    .B(net5215),
    .C(net5214),
    .Y(_00952_));
 INVx1_ASAP7_75t_R _06666_ (.A(_00952_),
    .Y(_00953_));
 NOR2x1_ASAP7_75t_R _06667_ (.A(_00328_),
    .B(_00953_),
    .Y(_00954_));
 OA21x2_ASAP7_75t_R _06668_ (.A1(_00948_),
    .A2(_00954_),
    .B(net5363),
    .Y(_00012_));
 INVx1_ASAP7_75t_R _06669_ (.A(_00316_),
    .Y(_00955_));
 INVx2_ASAP7_75t_R _06670_ (.A(net5201),
    .Y(_00956_));
 BUFx3_ASAP7_75t_R place3045 (.A(_05145_),
    .Y(net3045));
 AND3x1_ASAP7_75t_R _06672_ (.A(net5042),
    .B(net5041),
    .C(net5363),
    .Y(_00005_));
 INVx1_ASAP7_75t_R _06673_ (.A(_00069_),
    .Y(\tx_fifo.write_ptr[0] ));
 INVx1_ASAP7_75t_R _06674_ (.A(net5357),
    .Y(\tx_fifo.read_ptr[0] ));
 INVx1_ASAP7_75t_R _06675_ (.A(_00308_),
    .Y(\tx_fifo.write_ptr[1] ));
 INVx1_ASAP7_75t_R _06676_ (.A(net5356),
    .Y(\tx_fifo.read_ptr[1] ));
 NOR2x1_ASAP7_75t_R _06677_ (.A(_06525_),
    .B(_00316_),
    .Y(_00958_));
 BUFx3_ASAP7_75t_R place3043 (.A(_06233_),
    .Y(net3043));
 XOR2x2_ASAP7_75t_R _06679_ (.A(_00302_),
    .B(_00309_),
    .Y(_00960_));
 BUFx6f_ASAP7_75t_R place3042 (.A(_06241_),
    .Y(net3042));
 XOR2x2_ASAP7_75t_R _06681_ (.A(_00303_),
    .B(_00310_),
    .Y(_00962_));
 NOR2x1_ASAP7_75t_R _06682_ (.A(_00960_),
    .B(_00962_),
    .Y(_00963_));
 XNOR2x2_ASAP7_75t_R _06683_ (.A(_00304_),
    .B(_00311_),
    .Y(_00964_));
 XNOR2x2_ASAP7_75t_R _06684_ (.A(_00305_),
    .B(_00312_),
    .Y(_00965_));
 AND3x1_ASAP7_75t_R _06685_ (.A(_00963_),
    .B(_00964_),
    .C(_00965_),
    .Y(_00966_));
 XNOR2x2_ASAP7_75t_R _06686_ (.A(net5346),
    .B(_00313_),
    .Y(_00967_));
 XNOR2x2_ASAP7_75t_R _06687_ (.A(net5348),
    .B(_00544_),
    .Y(_00968_));
 XNOR2x2_ASAP7_75t_R _06688_ (.A(net5347),
    .B(_00314_),
    .Y(_00969_));
 XNOR2x2_ASAP7_75t_R _06689_ (.A(net5349),
    .B(_00543_),
    .Y(_00970_));
 AND4x1_ASAP7_75t_R _06690_ (.A(_00967_),
    .B(_00968_),
    .C(_00969_),
    .D(_00970_),
    .Y(_00971_));
 AND2x2_ASAP7_75t_R _06691_ (.A(_00966_),
    .B(_00971_),
    .Y(_00972_));
 INVx1_ASAP7_75t_R _06692_ (.A(_00972_),
    .Y(_00973_));
 AND2x2_ASAP7_75t_R _06693_ (.A(_00123_),
    .B(_00122_),
    .Y(_00974_));
 AND3x1_ASAP7_75t_R _06694_ (.A(_00974_),
    .B(_00120_),
    .C(_00121_),
    .Y(_00975_));
 AND2x2_ASAP7_75t_R _06695_ (.A(_00127_),
    .B(_00126_),
    .Y(_00976_));
 AND3x1_ASAP7_75t_R _06696_ (.A(_00976_),
    .B(_00124_),
    .C(_00125_),
    .Y(_00977_));
 AND2x2_ASAP7_75t_R _06697_ (.A(_00977_),
    .B(_00975_),
    .Y(_00978_));
 AND2x2_ASAP7_75t_R _06698_ (.A(_00118_),
    .B(_00119_),
    .Y(_00979_));
 AND3x1_ASAP7_75t_R _06699_ (.A(_00979_),
    .B(_00116_),
    .C(_00117_),
    .Y(_00980_));
 AND2x2_ASAP7_75t_R _06700_ (.A(_00112_),
    .B(_00114_),
    .Y(_00981_));
 AND5x1_ASAP7_75t_R _06701_ (.A(_00111_),
    .B(_00978_),
    .C(_00115_),
    .D(_00980_),
    .E(_00981_),
    .Y(_00982_));
 AND2x2_ASAP7_75t_R _06702_ (.A(_00129_),
    .B(_00128_),
    .Y(_00983_));
 AND3x1_ASAP7_75t_R _06703_ (.A(_00983_),
    .B(net5168),
    .C(net5169),
    .Y(_00984_));
 AND2x2_ASAP7_75t_R _06704_ (.A(_00132_),
    .B(_00133_),
    .Y(_00985_));
 AND4x1_ASAP7_75t_R _06705_ (.A(_00984_),
    .B(net5146),
    .C(net5145),
    .D(net5035),
    .Y(_00986_));
 AND2x2_ASAP7_75t_R _06706_ (.A(_00106_),
    .B(_00107_),
    .Y(_00987_));
 AND3x1_ASAP7_75t_R _06707_ (.A(net5034),
    .B(net5149),
    .C(net5150),
    .Y(_00988_));
 INVx1_ASAP7_75t_R _06708_ (.A(_00110_),
    .Y(_00989_));
 INVx1_ASAP7_75t_R _06709_ (.A(net5153),
    .Y(_00990_));
 OR3x1_ASAP7_75t_R _06710_ (.A(_00536_),
    .B(_00990_),
    .C(_00989_),
    .Y(_00991_));
 INVx1_ASAP7_75t_R _06711_ (.A(_00991_),
    .Y(_00992_));
 AND2x4_ASAP7_75t_R _06712_ (.A(_00988_),
    .B(_00992_),
    .Y(_00993_));
 AND3x1_ASAP7_75t_R _06713_ (.A(net4697),
    .B(_00986_),
    .C(_00982_),
    .Y(_00994_));
 BUFx3_ASAP7_75t_R place3041 (.A(_06244_),
    .Y(net3041));
 OA21x2_ASAP7_75t_R _06715_ (.A1(_00994_),
    .A2(net5199),
    .B(_00162_),
    .Y(_00996_));
 NOR2x1_ASAP7_75t_R _06716_ (.A(_00973_),
    .B(_00996_),
    .Y(_00997_));
 INVx1_ASAP7_75t_R _06717_ (.A(_00997_),
    .Y(_00998_));
 BUFx3_ASAP7_75t_R place3040 (.A(_02193_),
    .Y(net3040));
 AND2x4_ASAP7_75t_R _06719_ (.A(net5202),
    .B(net5198),
    .Y(_01000_));
 AND2x4_ASAP7_75t_R _06720_ (.A(_00998_),
    .B(_01000_),
    .Y(_01001_));
 NOR2x1p5_ASAP7_75t_R _06721_ (.A(_06525_),
    .B(net4432),
    .Y(_00020_));
 AO21x1_ASAP7_75t_R _06722_ (.A1(net5041),
    .A2(_00958_),
    .B(_00020_),
    .Y(_00022_));
 NAND2x1p5_ASAP7_75t_R _06723_ (.A(net4432),
    .B(net5363),
    .Y(_00021_));
 INVx2_ASAP7_75t_R _06724_ (.A(net4577),
    .Y(_01002_));
 AND3x1_ASAP7_75t_R _06725_ (.A(_01002_),
    .B(net5363),
    .C(net4641),
    .Y(_00019_));
 INVx2_ASAP7_75t_R _06726_ (.A(net5199),
    .Y(_01003_));
 NOR2x1_ASAP7_75t_R _06727_ (.A(_00335_),
    .B(_00955_),
    .Y(_01004_));
 AO21x1_ASAP7_75t_R _06728_ (.A1(net4640),
    .A2(net5022),
    .B(net4855),
    .Y(_01005_));
 AND2x2_ASAP7_75t_R _06729_ (.A(_01005_),
    .B(net5363),
    .Y(_00018_));
 OA21x2_ASAP7_75t_R _06730_ (.A1(_00322_),
    .A2(_00330_),
    .B(net5204),
    .Y(_01006_));
 NOR2x1_ASAP7_75t_R _06731_ (.A(_01006_),
    .B(_00914_),
    .Y(_00016_));
 INVx1_ASAP7_75t_R _06732_ (.A(_00327_),
    .Y(_01007_));
 AO21x1_ASAP7_75t_R _06733_ (.A1(_01007_),
    .A2(_00072_),
    .B(net5360),
    .Y(_01008_));
 INVx1_ASAP7_75t_R _06734_ (.A(_01008_),
    .Y(_01009_));
 NAND2x1_ASAP7_75t_R _06735_ (.A(_00176_),
    .B(_01009_),
    .Y(_00011_));
 INVx2_ASAP7_75t_R _06736_ (.A(_00872_),
    .Y(\u_window_buffer.write_ptr[0] ));
 BUFx3_ASAP7_75t_R place3044 (.A(_06217_),
    .Y(net3044));
 BUFx3_ASAP7_75t_R place3039 (.A(_03907_),
    .Y(net3039));
 NOR2x2_ASAP7_75t_R _06739_ (.A(_00410_),
    .B(net4806),
    .Y(_01012_));
 BUFx3_ASAP7_75t_R place3038 (.A(_03917_),
    .Y(net3038));
 NOR2x2_ASAP7_75t_R _06741_ (.A(net4802),
    .B(net4804),
    .Y(_01014_));
 NAND2x1p5_ASAP7_75t_R _06742_ (.A(_01014_),
    .B(_01012_),
    .Y(_01015_));
 BUFx3_ASAP7_75t_R place3037 (.A(_05128_),
    .Y(net3037));
 NOR2x2_ASAP7_75t_R _06744_ (.A(net4797),
    .B(net4799),
    .Y(_01017_));
 BUFx3_ASAP7_75t_R place3036 (.A(_05136_),
    .Y(net3036));
 NOR2x2_ASAP7_75t_R _06746_ (.A(net4795),
    .B(net4793),
    .Y(_01019_));
 NAND2x1p5_ASAP7_75t_R _06747_ (.A(_01017_),
    .B(_01019_),
    .Y(_01020_));
 NOR2x1p5_ASAP7_75t_R _06748_ (.A(_01015_),
    .B(_01020_),
    .Y(_01021_));
 NOR2x2_ASAP7_75t_R _06749_ (.A(net4789),
    .B(net4791),
    .Y(_01022_));
 BUFx3_ASAP7_75t_R place3035 (.A(_05153_),
    .Y(net3035));
 NOR2x2_ASAP7_75t_R _06751_ (.A(net4787),
    .B(net4785),
    .Y(_01024_));
 NAND2x2_ASAP7_75t_R _06752_ (.A(_01022_),
    .B(_01024_),
    .Y(_01025_));
 BUFx3_ASAP7_75t_R place3034 (.A(_05161_),
    .Y(net3034));
 NOR2x2_ASAP7_75t_R _06754_ (.A(net4781),
    .B(net4783),
    .Y(_01027_));
 OAI21x1_ASAP7_75t_R _06755_ (.A1(net4830),
    .A2(net4779),
    .B(_00437_),
    .Y(_01028_));
 OAI21x1_ASAP7_75t_R _06756_ (.A1(_00435_),
    .A2(net4783),
    .B(_00433_),
    .Y(_01029_));
 AOI21x1_ASAP7_75t_R _06757_ (.A1(_01027_),
    .A2(_01028_),
    .B(_01029_),
    .Y(_01030_));
 OAI21x1_ASAP7_75t_R _06758_ (.A1(_00431_),
    .A2(net4787),
    .B(_00429_),
    .Y(_01031_));
 OAI21x1_ASAP7_75t_R _06759_ (.A1(net4831),
    .A2(net4791),
    .B(_00425_),
    .Y(_01032_));
 AOI21x1_ASAP7_75t_R _06760_ (.A1(_01022_),
    .A2(_01031_),
    .B(_01032_),
    .Y(_01033_));
 OAI21x1_ASAP7_75t_R _06761_ (.A1(_01025_),
    .A2(_01030_),
    .B(_01033_),
    .Y(_01034_));
 OAI21x1_ASAP7_75t_R _06762_ (.A1(_00423_),
    .A2(net4795),
    .B(_00421_),
    .Y(_01035_));
 OAI21x1_ASAP7_75t_R _06763_ (.A1(_00419_),
    .A2(net4800),
    .B(_00417_),
    .Y(_01036_));
 AOI21x1_ASAP7_75t_R _06764_ (.A1(_01017_),
    .A2(_01035_),
    .B(_01036_),
    .Y(_01037_));
 OAI21x1_ASAP7_75t_R _06765_ (.A1(net4832),
    .A2(net4805),
    .B(_00413_),
    .Y(_01038_));
 OAI21x1_ASAP7_75t_R _06766_ (.A1(_00411_),
    .A2(net4808),
    .B(_00409_),
    .Y(_01039_));
 AOI21x1_ASAP7_75t_R _06767_ (.A1(_01012_),
    .A2(_01038_),
    .B(_01039_),
    .Y(_01040_));
 OAI21x1_ASAP7_75t_R _06768_ (.A1(_01015_),
    .A2(_01037_),
    .B(_01040_),
    .Y(_01041_));
 AOI21x1_ASAP7_75t_R _06769_ (.A1(_01021_),
    .A2(_01034_),
    .B(_01041_),
    .Y(_01042_));
 NOR2x2_ASAP7_75t_R _06770_ (.A(net4766),
    .B(net4767),
    .Y(_01043_));
 NOR2x1_ASAP7_75t_R _06771_ (.A(net4765),
    .B(net4763),
    .Y(_01044_));
 NAND2x2_ASAP7_75t_R _06772_ (.A(_01043_),
    .B(_01044_),
    .Y(_01045_));
 NOR2x2_ASAP7_75t_R _06773_ (.A(net4773),
    .B(net4775),
    .Y(_01046_));
 NOR2x2_ASAP7_75t_R _06774_ (.A(net4769),
    .B(net4771),
    .Y(_01047_));
 NAND2x2_ASAP7_75t_R _06775_ (.A(_01047_),
    .B(_01046_),
    .Y(_01048_));
 OAI21x1_ASAP7_75t_R _06776_ (.A1(_00459_),
    .A2(net5364),
    .B(_00457_),
    .Y(_01049_));
 INVx1_ASAP7_75t_R _06777_ (.A(_01049_),
    .Y(_01050_));
 NOR3x2_ASAP7_75t_R _06778_ (.B(_01048_),
    .C(_01045_),
    .Y(_01051_),
    .A(_01050_));
 OAI21x1_ASAP7_75t_R _06779_ (.A1(net4825),
    .A2(net4765),
    .B(_00453_),
    .Y(_01052_));
 OAI21x1_ASAP7_75t_R _06780_ (.A1(net4767),
    .A2(_00451_),
    .B(_00449_),
    .Y(_01053_));
 AOI21x1_ASAP7_75t_R _06781_ (.A1(_01043_),
    .A2(net4714),
    .B(_01053_),
    .Y(_01054_));
 OAI21x1_ASAP7_75t_R _06782_ (.A1(_00447_),
    .A2(net4771),
    .B(_00445_),
    .Y(_01055_));
 OAI21x1_ASAP7_75t_R _06783_ (.A1(net4829),
    .A2(net4775),
    .B(_00441_),
    .Y(_01056_));
 AOI21x1_ASAP7_75t_R _06784_ (.A1(_01046_),
    .A2(_01055_),
    .B(_01056_),
    .Y(_01057_));
 OAI21x1_ASAP7_75t_R _06785_ (.A1(_01048_),
    .A2(_01054_),
    .B(_01057_),
    .Y(_01058_));
 BUFx3_ASAP7_75t_R place3033 (.A(_05164_),
    .Y(net3033));
 NOR2x2_ASAP7_75t_R _06787_ (.A(net4777),
    .B(net4779),
    .Y(_01060_));
 NAND2x2_ASAP7_75t_R _06788_ (.A(_01060_),
    .B(_01027_),
    .Y(_01061_));
 NOR2x2_ASAP7_75t_R _06789_ (.A(_01025_),
    .B(_01061_),
    .Y(_01062_));
 AND2x4_ASAP7_75t_R _06790_ (.A(_01062_),
    .B(_01021_),
    .Y(_01063_));
 OAI21x1_ASAP7_75t_R _06791_ (.A1(net5371),
    .A2(net5377),
    .B(_01063_),
    .Y(_01064_));
 NAND2x1_ASAP7_75t_R _06792_ (.A(_01042_),
    .B(_01064_),
    .Y(_01065_));
 BUFx3_ASAP7_75t_R place3032 (.A(_05178_),
    .Y(net3032));
 NOR2x1_ASAP7_75t_R _06794_ (.A(_00406_),
    .B(net5375),
    .Y(_01067_));
 INVx1_ASAP7_75t_R _06795_ (.A(_00404_),
    .Y(_01068_));
 INVx1_ASAP7_75t_R _06796_ (.A(_00402_),
    .Y(_01069_));
 AND3x1_ASAP7_75t_R _06797_ (.A(net4713),
    .B(_01068_),
    .C(_01069_),
    .Y(_01070_));
 OA21x2_ASAP7_75t_R _06798_ (.A1(_00407_),
    .A2(net4812),
    .B(_00405_),
    .Y(_01071_));
 OA21x2_ASAP7_75t_R _06799_ (.A1(_01071_),
    .A2(_00404_),
    .B(_00403_),
    .Y(_01072_));
 OAI21x1_ASAP7_75t_R _06800_ (.A1(_00402_),
    .A2(_01072_),
    .B(_00401_),
    .Y(_01073_));
 AO21x1_ASAP7_75t_R _06801_ (.A1(_01065_),
    .A2(_01070_),
    .B(_01073_),
    .Y(_01074_));
 XNOR2x2_ASAP7_75t_R _06802_ (.A(_00080_),
    .B(_00139_),
    .Y(_01075_));
 XOR2x2_ASAP7_75t_R _06803_ (.A(_01074_),
    .B(_01075_),
    .Y(_01076_));
 INVx2_ASAP7_75t_R _06804_ (.A(_01076_),
    .Y(_01077_));
 BUFx3_ASAP7_75t_R place3031 (.A(_06245_),
    .Y(net3031));
 BUFx3_ASAP7_75t_R place3030 (.A(net5458),
    .Y(net3030));
 INVx1_ASAP7_75t_R _06807_ (.A(net4761),
    .Y(_01080_));
 NOR2x1_ASAP7_75t_R _06808_ (.A(_01080_),
    .B(net4287),
    .Y(_01081_));
 AO21x1_ASAP7_75t_R _06809_ (.A1(net4658),
    .A2(net4287),
    .B(_01081_),
    .Y(_00465_));
 INVx2_ASAP7_75t_R _06810_ (.A(_00071_),
    .Y(\u_window_buffer.write_ptr[1] ));
 BUFx3_ASAP7_75t_R place3029 (.A(_02210_),
    .Y(net3029));
 INVx5_ASAP7_75t_R _06812_ (.A(_00461_),
    .Y(\u_window_buffer.read_ptr[0] ));
 BUFx3_ASAP7_75t_R place3028 (.A(_02218_),
    .Y(net3028));
 OA21x2_ASAP7_75t_R _06814_ (.A1(_00343_),
    .A2(_00345_),
    .B(_00342_),
    .Y(_01084_));
 OAI21x1_ASAP7_75t_R _06815_ (.A1(net4644),
    .A2(_00357_),
    .B(_00354_),
    .Y(_01085_));
 AND2x2_ASAP7_75t_R _06816_ (.A(_00227_),
    .B(net5281),
    .Y(_01086_));
 OA21x2_ASAP7_75t_R _06817_ (.A1(_01086_),
    .A2(_00371_),
    .B(_00370_),
    .Y(_01087_));
 OA21x2_ASAP7_75t_R _06818_ (.A1(_01087_),
    .A2(_00364_),
    .B(_00363_),
    .Y(_01088_));
 OAI21x1_ASAP7_75t_R _06819_ (.A1(_00361_),
    .A2(_01088_),
    .B(_00360_),
    .Y(_01089_));
 INVx1_ASAP7_75t_R _06820_ (.A(_00355_),
    .Y(_01090_));
 INVx1_ASAP7_75t_R _06821_ (.A(_00358_),
    .Y(_01091_));
 AND3x1_ASAP7_75t_R _06822_ (.A(_01089_),
    .B(_01091_),
    .C(_01090_),
    .Y(_01092_));
 INVx1_ASAP7_75t_R _06823_ (.A(_00352_),
    .Y(_01093_));
 OAI21x1_ASAP7_75t_R _06824_ (.A1(_01085_),
    .A2(_01092_),
    .B(_01093_),
    .Y(_01094_));
 AO21x1_ASAP7_75t_R _06825_ (.A1(_01094_),
    .A2(_00351_),
    .B(_00349_),
    .Y(_01095_));
 OR2x2_ASAP7_75t_R _06826_ (.A(_00343_),
    .B(_00346_),
    .Y(_01096_));
 AO21x1_ASAP7_75t_R _06827_ (.A1(_01095_),
    .A2(_00348_),
    .B(_01096_),
    .Y(_01097_));
 AO32x1_ASAP7_75t_R _06828_ (.A1(_00236_),
    .A2(_00873_),
    .A3(_00879_),
    .B1(_01084_),
    .B2(_01097_),
    .Y(_01098_));
 INVx2_ASAP7_75t_R _06829_ (.A(_01098_),
    .Y(_01099_));
 NOR2x1p5_ASAP7_75t_R _06830_ (.A(net5329),
    .B(net4224),
    .Y(_01100_));
 AND2x2_ASAP7_75t_R _06831_ (.A(_00067_),
    .B(_00488_),
    .Y(_01101_));
 BUFx3_ASAP7_75t_R place3048 (.A(_03940_),
    .Y(net3048));
 AO32x1_ASAP7_75t_R _06833_ (.A1(_00481_),
    .A2(_01101_),
    .A3(_00480_),
    .B1(net5259),
    .B2(_00057_),
    .Y(_01103_));
 INVx1_ASAP7_75t_R _06834_ (.A(_00068_),
    .Y(_01104_));
 AND2x2_ASAP7_75t_R _06835_ (.A(_01103_),
    .B(_01104_),
    .Y(_01105_));
 INVx1_ASAP7_75t_R _06836_ (.A(_00389_),
    .Y(_01106_));
 INVx1_ASAP7_75t_R _06837_ (.A(_00495_),
    .Y(_01107_));
 OA21x2_ASAP7_75t_R _06838_ (.A1(_01107_),
    .A2(_00400_),
    .B(_00399_),
    .Y(_01108_));
 OA21x2_ASAP7_75t_R _06839_ (.A1(_01108_),
    .A2(_00395_),
    .B(_00394_),
    .Y(_01109_));
 OAI21x1_ASAP7_75t_R _06840_ (.A1(_00392_),
    .A2(_01109_),
    .B(_00391_),
    .Y(_01110_));
 NAND2x1_ASAP7_75t_R _06841_ (.A(_01106_),
    .B(_01110_),
    .Y(_01111_));
 AO21x1_ASAP7_75t_R _06842_ (.A1(_01111_),
    .A2(_00388_),
    .B(_00386_),
    .Y(_01112_));
 AO21x1_ASAP7_75t_R _06843_ (.A1(_01112_),
    .A2(_00385_),
    .B(_00383_),
    .Y(_01113_));
 AO21x1_ASAP7_75t_R _06844_ (.A1(_01113_),
    .A2(_00382_),
    .B(_00380_),
    .Y(_01114_));
 AOI211x1_ASAP7_75t_R _06845_ (.A1(_01114_),
    .A2(_00379_),
    .B(_00374_),
    .C(_00377_),
    .Y(_01115_));
 OAI21x1_ASAP7_75t_R _06846_ (.A1(_00374_),
    .A2(_00376_),
    .B(_00373_),
    .Y(_01116_));
 AO21x1_ASAP7_75t_R _06847_ (.A1(_00890_),
    .A2(net5266),
    .B(net5265),
    .Y(_01117_));
 OA21x2_ASAP7_75t_R _06848_ (.A1(_01116_),
    .A2(_01115_),
    .B(_01117_),
    .Y(_01118_));
 NOR2x1p5_ASAP7_75t_R _06849_ (.A(net5330),
    .B(net4235),
    .Y(_01119_));
 BUFx6f_ASAP7_75t_R place3026 (.A(_02226_),
    .Y(net3026));
 OR3x1_ASAP7_75t_R _06851_ (.A(net4152),
    .B(net4179),
    .C(_01105_),
    .Y(_01121_));
 NOR2x1_ASAP7_75t_R _06852_ (.A(net5332),
    .B(net5222),
    .Y(_01122_));
 OA21x2_ASAP7_75t_R _06853_ (.A1(_01121_),
    .A2(_01122_),
    .B(net211),
    .Y(_00010_));
 INVx2_ASAP7_75t_R _06854_ (.A(_00184_),
    .Y(_01123_));
 NOR2x1p5_ASAP7_75t_R _06855_ (.A(_00323_),
    .B(_01123_),
    .Y(_01124_));
 INVx1_ASAP7_75t_R _06856_ (.A(_00294_),
    .Y(_01125_));
 OR3x1_ASAP7_75t_R _06857_ (.A(_01124_),
    .B(net5361),
    .C(_01125_),
    .Y(_00008_));
 NOR2x1_ASAP7_75t_R _06858_ (.A(net5330),
    .B(net4854),
    .Y(_01126_));
 AND3x1_ASAP7_75t_R _06859_ (.A(net4235),
    .B(net4224),
    .C(net4747),
    .Y(_01127_));
 AND4x1_ASAP7_75t_R _06860_ (.A(_00246_),
    .B(_00247_),
    .C(_00248_),
    .D(_00249_),
    .Y(_01128_));
 INVx1_ASAP7_75t_R _06861_ (.A(_00245_),
    .Y(_01129_));
 AND3x1_ASAP7_75t_R _06862_ (.A(_01128_),
    .B(_00244_),
    .C(_01129_),
    .Y(_01130_));
 AND5x2_ASAP7_75t_R _06863_ (.A(_01130_),
    .B(_00250_),
    .C(_00251_),
    .D(_00252_),
    .E(_00253_),
    .Y(_01131_));
 NOR2x2_ASAP7_75t_R _06864_ (.A(net4746),
    .B(net5331),
    .Y(_01132_));
 BUFx3_ASAP7_75t_R place3025 (.A(_03913_),
    .Y(net3025));
 OA21x2_ASAP7_75t_R _06866_ (.A1(_01127_),
    .A2(net4696),
    .B(net5362),
    .Y(_00009_));
 AO32x1_ASAP7_75t_R _06867_ (.A1(net5022),
    .A2(_00316_),
    .A3(_00956_),
    .B1(net4641),
    .B2(_01002_),
    .Y(_01134_));
 AND3x4_ASAP7_75t_R _06868_ (.A(_00336_),
    .B(_00335_),
    .C(_00055_),
    .Y(_01135_));
 AND3x1_ASAP7_75t_R _06869_ (.A(net5016),
    .B(_00162_),
    .C(net5202),
    .Y(_01136_));
 NOR2x1_ASAP7_75t_R _06870_ (.A(net4855),
    .B(net4853),
    .Y(_01137_));
 OA21x2_ASAP7_75t_R _06871_ (.A1(_00054_),
    .A2(_01137_),
    .B(_01001_),
    .Y(_01138_));
 AND2x2_ASAP7_75t_R _06872_ (.A(_00056_),
    .B(_00316_),
    .Y(_01139_));
 INVx1_ASAP7_75t_R _06873_ (.A(_01136_),
    .Y(_01140_));
 OA21x2_ASAP7_75t_R _06874_ (.A1(net5201),
    .A2(_01139_),
    .B(_01140_),
    .Y(_01141_));
 AO32x1_ASAP7_75t_R _06875_ (.A1(_01000_),
    .A2(_00998_),
    .A3(_01141_),
    .B1(_00056_),
    .B2(net4853),
    .Y(_01142_));
 XNOR2x2_ASAP7_75t_R _06876_ (.A(_01138_),
    .B(_01142_),
    .Y(_01143_));
 XOR2x2_ASAP7_75t_R _06877_ (.A(net4762),
    .B(net4823),
    .Y(_01144_));
 INVx1_ASAP7_75t_R _06878_ (.A(_01144_),
    .Y(_01145_));
 AND3x1_ASAP7_75t_R _06879_ (.A(_01145_),
    .B(net5143),
    .C(net4761),
    .Y(_01146_));
 NAND2x1_ASAP7_75t_R _06880_ (.A(net4825),
    .B(_00457_),
    .Y(_01147_));
 NOR2x1_ASAP7_75t_R _06881_ (.A(net5365),
    .B(_00460_),
    .Y(_01148_));
 NAND2x1_ASAP7_75t_R _06882_ (.A(net4825),
    .B(net4763),
    .Y(_01149_));
 OAI21x1_ASAP7_75t_R _06883_ (.A1(_01148_),
    .A2(_01147_),
    .B(_01149_),
    .Y(_01150_));
 INVx1_ASAP7_75t_R _06884_ (.A(net5435),
    .Y(_01151_));
 XOR2x2_ASAP7_75t_R _06885_ (.A(net4656),
    .B(_01151_),
    .Y(_01152_));
 INVx1_ASAP7_75t_R _06886_ (.A(net4764),
    .Y(_01153_));
 XOR2x2_ASAP7_75t_R _06887_ (.A(net4716),
    .B(_01153_),
    .Y(_01154_));
 INVx1_ASAP7_75t_R _06888_ (.A(net4654),
    .Y(_01155_));
 AND3x1_ASAP7_75t_R _06889_ (.A(_01146_),
    .B(_01152_),
    .C(_01155_),
    .Y(_01156_));
 INVx1_ASAP7_75t_R _06890_ (.A(_01156_),
    .Y(_01157_));
 NAND2x1_ASAP7_75t_R _06891_ (.A(net4494),
    .B(net4287),
    .Y(_01158_));
 AOI21x1_ASAP7_75t_R _06892_ (.A1(_01049_),
    .A2(_01044_),
    .B(net5432),
    .Y(_01159_));
 INVx1_ASAP7_75t_R _06893_ (.A(net4766),
    .Y(_01160_));
 XOR2x2_ASAP7_75t_R _06894_ (.A(net4653),
    .B(_01160_),
    .Y(_01161_));
 XOR2x2_ASAP7_75t_R _06895_ (.A(_01158_),
    .B(net4595),
    .Y(_01162_));
 INVx1_ASAP7_75t_R _06896_ (.A(_01162_),
    .Y(_01163_));
 NOR2x2_ASAP7_75t_R _06897_ (.A(net4766),
    .B(net4765),
    .Y(_01164_));
 INVx1_ASAP7_75t_R _06898_ (.A(_01164_),
    .Y(_01165_));
 OAI21x1_ASAP7_75t_R _06899_ (.A1(net4766),
    .A2(net4827),
    .B(net4828),
    .Y(_01166_));
 INVx1_ASAP7_75t_R _06900_ (.A(_01166_),
    .Y(_01167_));
 OAI21x1_ASAP7_75t_R _06901_ (.A1(_01165_),
    .A2(_01150_),
    .B(_01167_),
    .Y(_01168_));
 XOR2x2_ASAP7_75t_R _06902_ (.A(_01168_),
    .B(net4768),
    .Y(_01169_));
 AND3x1_ASAP7_75t_R _06903_ (.A(_01156_),
    .B(net4595),
    .C(net4538),
    .Y(_01170_));
 INVx1_ASAP7_75t_R _06904_ (.A(_01170_),
    .Y(_01171_));
 NAND2x1_ASAP7_75t_R _06905_ (.A(net4448),
    .B(net4287),
    .Y(_01172_));
 NAND2x1_ASAP7_75t_R _06906_ (.A(_01044_),
    .B(_01049_),
    .Y(_01173_));
 NOR2x1_ASAP7_75t_R _06907_ (.A(_01053_),
    .B(net5432),
    .Y(_01174_));
 NOR2x1_ASAP7_75t_R _06908_ (.A(_01043_),
    .B(_01053_),
    .Y(_01175_));
 AOI21x1_ASAP7_75t_R _06909_ (.A1(_01174_),
    .A2(_01173_),
    .B(_01175_),
    .Y(_01176_));
 XOR2x2_ASAP7_75t_R _06910_ (.A(net4770),
    .B(_01176_),
    .Y(_01177_));
 XOR2x2_ASAP7_75t_R _06911_ (.A(_01172_),
    .B(net4537),
    .Y(_01178_));
 INVx1_ASAP7_75t_R _06912_ (.A(_01178_),
    .Y(_01179_));
 NOR2x2_ASAP7_75t_R _06913_ (.A(net4773),
    .B(net4771),
    .Y(_01180_));
 NOR2x2_ASAP7_75t_R _06914_ (.A(net4769),
    .B(net4767),
    .Y(_01181_));
 NAND2x2_ASAP7_75t_R _06915_ (.A(_01180_),
    .B(_01181_),
    .Y(_01182_));
 NOR2x2_ASAP7_75t_R _06916_ (.A(net4775),
    .B(net4777),
    .Y(_01183_));
 NOR2x2_ASAP7_75t_R _06917_ (.A(net4781),
    .B(net5367),
    .Y(_01184_));
 NAND2x2_ASAP7_75t_R _06918_ (.A(_01183_),
    .B(_01184_),
    .Y(_01185_));
 NOR2x1_ASAP7_75t_R _06919_ (.A(_01182_),
    .B(_01185_),
    .Y(_01186_));
 NOR2x2_ASAP7_75t_R _06920_ (.A(net4785),
    .B(net4783),
    .Y(_01187_));
 NOR2x2_ASAP7_75t_R _06921_ (.A(net4789),
    .B(net4787),
    .Y(_01188_));
 NAND2x2_ASAP7_75t_R _06922_ (.A(_01187_),
    .B(_01188_),
    .Y(_01189_));
 NOR2x2_ASAP7_75t_R _06923_ (.A(net4793),
    .B(net4791),
    .Y(_01190_));
 NOR2x2_ASAP7_75t_R _06924_ (.A(net4795),
    .B(net4797),
    .Y(_01191_));
 NAND2x2_ASAP7_75t_R _06925_ (.A(_01190_),
    .B(_01191_),
    .Y(_01192_));
 NOR2x1_ASAP7_75t_R _06926_ (.A(_01189_),
    .B(_01192_),
    .Y(_01193_));
 NAND3x1_ASAP7_75t_R _06927_ (.A(_01168_),
    .B(_01186_),
    .C(_01193_),
    .Y(_01194_));
 OAI21x1_ASAP7_75t_R _06928_ (.A1(net4769),
    .A2(_00449_),
    .B(_00447_),
    .Y(_01195_));
 OAI21x1_ASAP7_75t_R _06929_ (.A1(net4773),
    .A2(_00445_),
    .B(_00443_),
    .Y(_01196_));
 AOI21x1_ASAP7_75t_R _06930_ (.A1(_01180_),
    .A2(_01195_),
    .B(_01196_),
    .Y(_01197_));
 OAI21x1_ASAP7_75t_R _06931_ (.A1(net4777),
    .A2(_00441_),
    .B(net5378),
    .Y(_01198_));
 OAI21x1_ASAP7_75t_R _06932_ (.A1(net4781),
    .A2(_00437_),
    .B(_00435_),
    .Y(_01199_));
 AOI21x1_ASAP7_75t_R _06933_ (.A1(_01184_),
    .A2(_01198_),
    .B(_01199_),
    .Y(_01200_));
 OAI21x1_ASAP7_75t_R _06934_ (.A1(_01185_),
    .A2(_01197_),
    .B(_01200_),
    .Y(_01201_));
 OAI21x1_ASAP7_75t_R _06935_ (.A1(net4785),
    .A2(_00433_),
    .B(_00431_),
    .Y(_01202_));
 OAI21x1_ASAP7_75t_R _06936_ (.A1(net4789),
    .A2(_00429_),
    .B(_00427_),
    .Y(_01203_));
 AOI21x1_ASAP7_75t_R _06937_ (.A1(_01188_),
    .A2(_01202_),
    .B(_01203_),
    .Y(_01204_));
 OAI21x1_ASAP7_75t_R _06938_ (.A1(net4793),
    .A2(_00425_),
    .B(_00423_),
    .Y(_01205_));
 OAI21x1_ASAP7_75t_R _06939_ (.A1(_00421_),
    .A2(net4798),
    .B(_00419_),
    .Y(_01206_));
 AOI21x1_ASAP7_75t_R _06940_ (.A1(_01191_),
    .A2(_01205_),
    .B(_01206_),
    .Y(_01207_));
 OAI21x1_ASAP7_75t_R _06941_ (.A1(net4651),
    .A2(net4650),
    .B(_01207_),
    .Y(_01208_));
 AOI21x1_ASAP7_75t_R _06942_ (.A1(net4592),
    .A2(_01201_),
    .B(_01208_),
    .Y(_01209_));
 AO21x1_ASAP7_75t_R _06943_ (.A1(_01194_),
    .A2(_01209_),
    .B(net4801),
    .Y(_01210_));
 NAND3x1_ASAP7_75t_R _06944_ (.A(_01194_),
    .B(_01209_),
    .C(net4801),
    .Y(_01211_));
 NAND2x1_ASAP7_75t_R _06945_ (.A(net4493),
    .B(net4492),
    .Y(_01212_));
 NAND2x2_ASAP7_75t_R _06946_ (.A(_01187_),
    .B(_01184_),
    .Y(_01213_));
 NAND2x2_ASAP7_75t_R _06947_ (.A(_01190_),
    .B(_01188_),
    .Y(_01214_));
 NOR2x2_ASAP7_75t_R _06948_ (.A(_01213_),
    .B(_01214_),
    .Y(_01215_));
 NAND2x2_ASAP7_75t_R _06949_ (.A(_01180_),
    .B(_01183_),
    .Y(_01216_));
 AOI21x1_ASAP7_75t_R _06950_ (.A1(_01181_),
    .A2(_01166_),
    .B(_01195_),
    .Y(_01217_));
 AOI21x1_ASAP7_75t_R _06951_ (.A1(_01183_),
    .A2(_01196_),
    .B(_01198_),
    .Y(_01218_));
 OAI21x1_ASAP7_75t_R _06952_ (.A1(_01216_),
    .A2(_01217_),
    .B(_01218_),
    .Y(_01219_));
 AOI21x1_ASAP7_75t_R _06953_ (.A1(_01187_),
    .A2(_01199_),
    .B(_01202_),
    .Y(_01220_));
 AOI21x1_ASAP7_75t_R _06954_ (.A1(_01190_),
    .A2(_01203_),
    .B(_01205_),
    .Y(_01221_));
 OAI21x1_ASAP7_75t_R _06955_ (.A1(_01214_),
    .A2(_01220_),
    .B(_01221_),
    .Y(_01222_));
 AOI21x1_ASAP7_75t_R _06956_ (.A1(_01215_),
    .A2(_01219_),
    .B(_01222_),
    .Y(_01223_));
 NAND2x2_ASAP7_75t_R _06957_ (.A(_01181_),
    .B(_01164_),
    .Y(_01224_));
 NOR2x1_ASAP7_75t_R _06958_ (.A(_01224_),
    .B(_01216_),
    .Y(_01225_));
 INVx1_ASAP7_75t_R _06959_ (.A(net4655),
    .Y(_01226_));
 NAND3x1_ASAP7_75t_R _06960_ (.A(_01225_),
    .B(_01226_),
    .C(_01215_),
    .Y(_01227_));
 AO21x2_ASAP7_75t_R _06961_ (.A1(_01223_),
    .A2(_01227_),
    .B(net4796),
    .Y(_01228_));
 NAND3x2_ASAP7_75t_R _06962_ (.B(net4796),
    .C(_01227_),
    .Y(_01229_),
    .A(_01223_));
 NAND2x2_ASAP7_75t_R _06963_ (.A(_01024_),
    .B(_01027_),
    .Y(_01230_));
 NAND2x2_ASAP7_75t_R _06964_ (.A(_01022_),
    .B(_01019_),
    .Y(_01231_));
 NOR2x2_ASAP7_75t_R _06965_ (.A(_01230_),
    .B(_01231_),
    .Y(_01232_));
 NAND2x2_ASAP7_75t_R _06966_ (.A(_01060_),
    .B(_01046_),
    .Y(_01233_));
 AOI21x1_ASAP7_75t_R _06967_ (.A1(_01053_),
    .A2(_01047_),
    .B(_01055_),
    .Y(_01234_));
 AOI21x1_ASAP7_75t_R _06968_ (.A1(_01060_),
    .A2(_01056_),
    .B(_01028_),
    .Y(_01235_));
 OAI21x1_ASAP7_75t_R _06969_ (.A1(_01233_),
    .A2(_01234_),
    .B(_01235_),
    .Y(_01236_));
 AOI21x1_ASAP7_75t_R _06970_ (.A1(_01024_),
    .A2(_01029_),
    .B(_01031_),
    .Y(_01237_));
 AOI21x1_ASAP7_75t_R _06971_ (.A1(_01019_),
    .A2(_01032_),
    .B(_01035_),
    .Y(_01238_));
 OAI21x1_ASAP7_75t_R _06972_ (.A1(net5402),
    .A2(_01237_),
    .B(_01238_),
    .Y(_01239_));
 AOI21x1_ASAP7_75t_R _06973_ (.A1(_01236_),
    .A2(_01232_),
    .B(_01239_),
    .Y(_01240_));
 NAND2x2_ASAP7_75t_R _06974_ (.A(_01043_),
    .B(_01047_),
    .Y(_01241_));
 NOR2x2_ASAP7_75t_R _06975_ (.A(_01241_),
    .B(_01233_),
    .Y(_01242_));
 INVx2_ASAP7_75t_R _06976_ (.A(net5381),
    .Y(_01243_));
 NAND3x1_ASAP7_75t_R _06977_ (.A(_01242_),
    .B(_01243_),
    .C(_01232_),
    .Y(_01244_));
 AO21x2_ASAP7_75t_R _06978_ (.A1(_01240_),
    .A2(_01244_),
    .B(net4798),
    .Y(_01245_));
 NAND3x1_ASAP7_75t_R _06979_ (.A(_01240_),
    .B(_01244_),
    .C(net4798),
    .Y(_01246_));
 AOI22x1_ASAP7_75t_R _06980_ (.A1(_01228_),
    .A2(_01229_),
    .B1(_01246_),
    .B2(_01245_),
    .Y(_01247_));
 INVx1_ASAP7_75t_R _06981_ (.A(net4788),
    .Y(_01248_));
 OAI21x1_ASAP7_75t_R _06982_ (.A1(net4655),
    .A2(_01224_),
    .B(_01217_),
    .Y(_01249_));
 NOR2x1p5_ASAP7_75t_R _06983_ (.A(_01213_),
    .B(_01216_),
    .Y(_01250_));
 OAI21x1_ASAP7_75t_R _06984_ (.A1(_01213_),
    .A2(_01218_),
    .B(_01220_),
    .Y(_01251_));
 AO21x2_ASAP7_75t_R _06985_ (.A1(_01249_),
    .A2(net4588),
    .B(_01251_),
    .Y(_01252_));
 NOR2x1_ASAP7_75t_R _06986_ (.A(_01248_),
    .B(_01252_),
    .Y(_01253_));
 AND2x2_ASAP7_75t_R _06987_ (.A(_01252_),
    .B(_01248_),
    .Y(_01254_));
 NOR2x1_ASAP7_75t_R _06988_ (.A(_01230_),
    .B(_01233_),
    .Y(_01255_));
 OAI21x1_ASAP7_75t_R _06989_ (.A1(_01241_),
    .A2(_01159_),
    .B(_01234_),
    .Y(_01256_));
 OAI21x1_ASAP7_75t_R _06990_ (.A1(net5767),
    .A2(_01235_),
    .B(_01237_),
    .Y(_01257_));
 AOI21x1_ASAP7_75t_R _06991_ (.A1(net4587),
    .A2(_01256_),
    .B(_01257_),
    .Y(_01258_));
 XNOR2x2_ASAP7_75t_R _06992_ (.A(net4790),
    .B(_01258_),
    .Y(_01259_));
 OAI21x1_ASAP7_75t_R _06993_ (.A1(_01253_),
    .A2(_01254_),
    .B(_01259_),
    .Y(_01260_));
 INVx1_ASAP7_75t_R _06994_ (.A(net4445),
    .Y(_01261_));
 NOR2x2_ASAP7_75t_R _06995_ (.A(_01185_),
    .B(_01189_),
    .Y(_01262_));
 OAI21x1_ASAP7_75t_R _06996_ (.A1(net4764),
    .A2(net4824),
    .B(net4826),
    .Y(_01263_));
 AOI21x1_ASAP7_75t_R _06997_ (.A1(_01164_),
    .A2(_01263_),
    .B(_01166_),
    .Y(_01264_));
 OAI21x1_ASAP7_75t_R _06998_ (.A1(_01182_),
    .A2(_01264_),
    .B(_01197_),
    .Y(_01265_));
 OAI21x1_ASAP7_75t_R _06999_ (.A1(_01189_),
    .A2(_01200_),
    .B(_01204_),
    .Y(_01266_));
 AOI21x1_ASAP7_75t_R _07000_ (.A1(net4586),
    .A2(_01265_),
    .B(net4584),
    .Y(_01267_));
 NOR2x2_ASAP7_75t_R _07001_ (.A(net4764),
    .B(net4762),
    .Y(_01268_));
 NAND2x1_ASAP7_75t_R _07002_ (.A(_01164_),
    .B(_01268_),
    .Y(_01269_));
 NOR2x1_ASAP7_75t_R _07003_ (.A(_01269_),
    .B(net4652),
    .Y(_01270_));
 INVx1_ASAP7_75t_R _07004_ (.A(net4823),
    .Y(_01271_));
 NAND3x1_ASAP7_75t_R _07005_ (.A(_01270_),
    .B(net4585),
    .C(_01271_),
    .Y(_01272_));
 AO21x1_ASAP7_75t_R _07006_ (.A1(_01267_),
    .A2(_01272_),
    .B(net4792),
    .Y(_01273_));
 NAND3x1_ASAP7_75t_R _07007_ (.A(_01267_),
    .B(net4792),
    .C(_01272_),
    .Y(_01274_));
 AOI21x1_ASAP7_75t_R _07008_ (.A1(net4599),
    .A2(net5758),
    .B(_01034_),
    .Y(_01275_));
 NOR2x1_ASAP7_75t_R _07009_ (.A(_01045_),
    .B(net4657),
    .Y(_01276_));
 NAND3x1_ASAP7_75t_R _07010_ (.A(_01276_),
    .B(_01062_),
    .C(net4715),
    .Y(_01277_));
 AO21x2_ASAP7_75t_R _07011_ (.A1(_01275_),
    .A2(_01277_),
    .B(net4794),
    .Y(_01278_));
 NAND3x1_ASAP7_75t_R _07012_ (.A(_01275_),
    .B(_01277_),
    .C(net4794),
    .Y(_01279_));
 AOI22x1_ASAP7_75t_R _07013_ (.A1(_01273_),
    .A2(_01274_),
    .B1(_01278_),
    .B2(net5384),
    .Y(_01280_));
 NAND2x1_ASAP7_75t_R _07014_ (.A(_01261_),
    .B(_01280_),
    .Y(_01281_));
 INVx1_ASAP7_75t_R _07015_ (.A(net4782),
    .Y(_01282_));
 AOI211x1_ASAP7_75t_R _07016_ (.A1(_01243_),
    .A2(_01242_),
    .B(_01236_),
    .C(_01282_),
    .Y(_01283_));
 NAND2x1_ASAP7_75t_R _07017_ (.A(_01242_),
    .B(_01243_),
    .Y(_01284_));
 INVx2_ASAP7_75t_R _07018_ (.A(_01236_),
    .Y(_01285_));
 AOI21x1_ASAP7_75t_R _07019_ (.A1(_01285_),
    .A2(_01284_),
    .B(net4782),
    .Y(_01286_));
 NOR3x1_ASAP7_75t_R _07020_ (.A(net4655),
    .B(_01224_),
    .C(_01216_),
    .Y(_01287_));
 INVx1_ASAP7_75t_R _07021_ (.A(net4780),
    .Y(_01288_));
 NOR3x1_ASAP7_75t_R _07022_ (.A(_01287_),
    .B(_01219_),
    .C(_01288_),
    .Y(_01289_));
 INVx1_ASAP7_75t_R _07023_ (.A(_01219_),
    .Y(_01290_));
 INVx1_ASAP7_75t_R _07024_ (.A(_01287_),
    .Y(_01291_));
 AOI21x1_ASAP7_75t_R _07025_ (.A1(_01290_),
    .A2(_01291_),
    .B(net4780),
    .Y(_01292_));
 OAI22x1_ASAP7_75t_R _07026_ (.A1(_01283_),
    .A2(_01286_),
    .B1(_01289_),
    .B2(_01292_),
    .Y(_01293_));
 NOR2x1_ASAP7_75t_R _07027_ (.A(_01061_),
    .B(_01048_),
    .Y(_01294_));
 OAI21x1_ASAP7_75t_R _07028_ (.A1(_01061_),
    .A2(_01057_),
    .B(_01030_),
    .Y(_01295_));
 INVx1_ASAP7_75t_R _07029_ (.A(net4786),
    .Y(_01296_));
 AOI211x1_ASAP7_75t_R _07030_ (.A1(_01176_),
    .A2(_01294_),
    .B(_01295_),
    .C(_01296_),
    .Y(_01297_));
 INVx1_ASAP7_75t_R _07031_ (.A(_01295_),
    .Y(_01298_));
 NAND2x1_ASAP7_75t_R _07032_ (.A(_01294_),
    .B(_01176_),
    .Y(_01299_));
 AOI21x1_ASAP7_75t_R _07033_ (.A1(_01298_),
    .A2(_01299_),
    .B(net4786),
    .Y(_01300_));
 INVx1_ASAP7_75t_R _07034_ (.A(net4784),
    .Y(_01301_));
 AOI211x1_ASAP7_75t_R _07035_ (.A1(_01168_),
    .A2(net4593),
    .B(_01201_),
    .C(_01301_),
    .Y(_01302_));
 INVx1_ASAP7_75t_R _07036_ (.A(_01201_),
    .Y(_01303_));
 NAND2x1_ASAP7_75t_R _07037_ (.A(net4593),
    .B(net4594),
    .Y(_01304_));
 AOI21x1_ASAP7_75t_R _07038_ (.A1(_01303_),
    .A2(_01304_),
    .B(net4784),
    .Y(_01305_));
 OAI22x1_ASAP7_75t_R _07039_ (.A1(_01297_),
    .A2(_01300_),
    .B1(_01302_),
    .B2(_01305_),
    .Y(_01306_));
 NOR2x1_ASAP7_75t_R _07040_ (.A(_01293_),
    .B(_01306_),
    .Y(_01307_));
 XOR2x2_ASAP7_75t_R _07041_ (.A(_01249_),
    .B(net4772),
    .Y(_01308_));
 XOR2x2_ASAP7_75t_R _07042_ (.A(_01256_),
    .B(net4774),
    .Y(_01309_));
 NAND2x1_ASAP7_75t_R _07043_ (.A(_01308_),
    .B(_01309_),
    .Y(_01310_));
 NOR3x1_ASAP7_75t_R _07044_ (.A(_01269_),
    .B(_01182_),
    .C(net4823),
    .Y(_01311_));
 INVx1_ASAP7_75t_R _07045_ (.A(net4776),
    .Y(_01312_));
 NOR3x1_ASAP7_75t_R _07046_ (.A(net5404),
    .B(_01265_),
    .C(_01312_),
    .Y(_01313_));
 INVx1_ASAP7_75t_R _07047_ (.A(_01265_),
    .Y(_01314_));
 INVx1_ASAP7_75t_R _07048_ (.A(_01311_),
    .Y(_01315_));
 AOI21x1_ASAP7_75t_R _07049_ (.A1(_01314_),
    .A2(_01315_),
    .B(net4776),
    .Y(_01316_));
 INVx1_ASAP7_75t_R _07050_ (.A(net4778),
    .Y(_01317_));
 NOR3x1_ASAP7_75t_R _07051_ (.A(_01051_),
    .B(_01317_),
    .C(_01058_),
    .Y(_01318_));
 INVx1_ASAP7_75t_R _07052_ (.A(_01058_),
    .Y(_01319_));
 INVx1_ASAP7_75t_R _07053_ (.A(_01051_),
    .Y(_01320_));
 AOI21x1_ASAP7_75t_R _07054_ (.A1(_01319_),
    .A2(_01320_),
    .B(net4778),
    .Y(_01321_));
 OAI22x1_ASAP7_75t_R _07055_ (.A1(_01313_),
    .A2(_01316_),
    .B1(net5370),
    .B2(_01321_),
    .Y(_01322_));
 NOR2x1_ASAP7_75t_R _07056_ (.A(_01322_),
    .B(_01310_),
    .Y(_01323_));
 NAND2x1_ASAP7_75t_R _07057_ (.A(_01169_),
    .B(_01177_),
    .Y(_01324_));
 OR3x1_ASAP7_75t_R _07058_ (.A(_01154_),
    .B(_00463_),
    .C(_01144_),
    .Y(_01325_));
 INVx1_ASAP7_75t_R _07059_ (.A(_01325_),
    .Y(_01326_));
 NAND3x2_ASAP7_75t_R _07060_ (.B(_01161_),
    .C(_01152_),
    .Y(_01327_),
    .A(_01326_));
 NOR2x1_ASAP7_75t_R _07061_ (.A(_01324_),
    .B(_01327_),
    .Y(_01328_));
 NAND3x1_ASAP7_75t_R _07062_ (.A(_01307_),
    .B(_01323_),
    .C(_01328_),
    .Y(_01329_));
 NOR2x1_ASAP7_75t_R _07063_ (.A(net4339),
    .B(net4338),
    .Y(_01330_));
 BUFx3_ASAP7_75t_R place3024 (.A(_03918_),
    .Y(net3024));
 AOI21x1_ASAP7_75t_R _07065_ (.A1(net4447),
    .A2(_01330_),
    .B(net4341),
    .Y(_01332_));
 XNOR2x2_ASAP7_75t_R _07066_ (.A(_01212_),
    .B(_01332_),
    .Y(_01333_));
 INVx1_ASAP7_75t_R _07067_ (.A(net4176),
    .Y(_01334_));
 AOI22x1_ASAP7_75t_R _07068_ (.A1(_01210_),
    .A2(_01211_),
    .B1(_01246_),
    .B2(_01245_),
    .Y(_01335_));
 NOR2x1_ASAP7_75t_R _07069_ (.A(_01020_),
    .B(_01025_),
    .Y(_01336_));
 NAND3x1_ASAP7_75t_R _07070_ (.A(_01336_),
    .B(_01294_),
    .C(_01176_),
    .Y(_01337_));
 OAI21x1_ASAP7_75t_R _07071_ (.A1(_01020_),
    .A2(_01033_),
    .B(_01037_),
    .Y(_01338_));
 AOI21x1_ASAP7_75t_R _07072_ (.A1(_01336_),
    .A2(_01295_),
    .B(_01338_),
    .Y(_01339_));
 NAND3x1_ASAP7_75t_R _07073_ (.A(net4803),
    .B(_01339_),
    .C(_01337_),
    .Y(_01340_));
 AO21x2_ASAP7_75t_R _07074_ (.A1(_01337_),
    .A2(_01339_),
    .B(net4803),
    .Y(_01341_));
 NOR2x2_ASAP7_75t_R _07075_ (.A(net5369),
    .B(net5366),
    .Y(_01342_));
 NAND2x1p5_ASAP7_75t_R _07076_ (.A(_01342_),
    .B(_01191_),
    .Y(_01343_));
 NOR2x1_ASAP7_75t_R _07077_ (.A(_01214_),
    .B(_01343_),
    .Y(_01344_));
 AND2x2_ASAP7_75t_R _07078_ (.A(_01250_),
    .B(_01344_),
    .Y(_01345_));
 NAND2x2_ASAP7_75t_R _07079_ (.A(_01249_),
    .B(_01345_),
    .Y(_01346_));
 OAI21x1_ASAP7_75t_R _07080_ (.A1(net4802),
    .A2(_00417_),
    .B(_00415_),
    .Y(_01347_));
 AOI21x1_ASAP7_75t_R _07081_ (.A1(_01342_),
    .A2(_01206_),
    .B(_01347_),
    .Y(_01348_));
 OAI21x1_ASAP7_75t_R _07082_ (.A1(net4649),
    .A2(_01221_),
    .B(_01348_),
    .Y(_01349_));
 AOI21x1_ASAP7_75t_R _07083_ (.A1(_01344_),
    .A2(_01251_),
    .B(_01349_),
    .Y(_01350_));
 NAND3x1_ASAP7_75t_R _07084_ (.A(_01346_),
    .B(_01350_),
    .C(net4805),
    .Y(_01351_));
 INVx1_ASAP7_75t_R _07085_ (.A(_01350_),
    .Y(_01352_));
 INVx2_ASAP7_75t_R _07086_ (.A(_01346_),
    .Y(_01353_));
 INVx1_ASAP7_75t_R _07087_ (.A(net4805),
    .Y(_01354_));
 OAI21x1_ASAP7_75t_R _07088_ (.A1(_01352_),
    .A2(_01353_),
    .B(_01354_),
    .Y(_01355_));
 AOI22x1_ASAP7_75t_R _07089_ (.A1(_01340_),
    .A2(_01341_),
    .B1(_01351_),
    .B2(_01355_),
    .Y(_01356_));
 NAND2x1_ASAP7_75t_R _07090_ (.A(_01356_),
    .B(_01335_),
    .Y(_01357_));
 NOR2x2_ASAP7_75t_R _07091_ (.A(net4804),
    .B(net4806),
    .Y(_01358_));
 NAND2x1_ASAP7_75t_R _07092_ (.A(_01342_),
    .B(_01358_),
    .Y(_01359_));
 NOR2x1_ASAP7_75t_R _07093_ (.A(_01192_),
    .B(_01359_),
    .Y(_01360_));
 AND2x2_ASAP7_75t_R _07094_ (.A(_01262_),
    .B(_01360_),
    .Y(_01361_));
 OAI21x1_ASAP7_75t_R _07095_ (.A1(net5403),
    .A2(_01265_),
    .B(_01361_),
    .Y(_01362_));
 OAI21x1_ASAP7_75t_R _07096_ (.A1(net4807),
    .A2(_00413_),
    .B(_00411_),
    .Y(_01363_));
 AOI21x1_ASAP7_75t_R _07097_ (.A1(net4710),
    .A2(_01347_),
    .B(_01363_),
    .Y(_01364_));
 OAI21x1_ASAP7_75t_R _07098_ (.A1(_01359_),
    .A2(_01207_),
    .B(_01364_),
    .Y(_01365_));
 AOI21x1_ASAP7_75t_R _07099_ (.A1(_01360_),
    .A2(_01266_),
    .B(_01365_),
    .Y(_01366_));
 NAND3x1_ASAP7_75t_R _07100_ (.A(net4809),
    .B(_01362_),
    .C(_01366_),
    .Y(_01367_));
 INVx1_ASAP7_75t_R _07101_ (.A(_01366_),
    .Y(_01368_));
 NAND2x1_ASAP7_75t_R _07102_ (.A(net4586),
    .B(net4581),
    .Y(_01369_));
 AOI21x1_ASAP7_75t_R _07103_ (.A1(_01314_),
    .A2(_01315_),
    .B(_01369_),
    .Y(_01370_));
 INVx1_ASAP7_75t_R _07104_ (.A(net4809),
    .Y(_01371_));
 OAI21x1_ASAP7_75t_R _07105_ (.A1(_01368_),
    .A2(_01370_),
    .B(_01371_),
    .Y(_01372_));
 NAND2x1p5_ASAP7_75t_R _07106_ (.A(_01014_),
    .B(_01017_),
    .Y(_01373_));
 NOR2x1_ASAP7_75t_R _07107_ (.A(_01231_),
    .B(_01373_),
    .Y(_01374_));
 AND2x2_ASAP7_75t_R _07108_ (.A(_01255_),
    .B(_01374_),
    .Y(_01375_));
 NAND2x1_ASAP7_75t_R _07109_ (.A(_01375_),
    .B(_01256_),
    .Y(_01376_));
 AOI21x1_ASAP7_75t_R _07110_ (.A1(net4717),
    .A2(_01036_),
    .B(_01038_),
    .Y(_01377_));
 OAI21x1_ASAP7_75t_R _07111_ (.A1(net4647),
    .A2(_01238_),
    .B(_01377_),
    .Y(_01378_));
 AOI21x1_ASAP7_75t_R _07112_ (.A1(net4580),
    .A2(_01257_),
    .B(_01378_),
    .Y(_01379_));
 AO21x2_ASAP7_75t_R _07113_ (.A1(_01376_),
    .A2(_01379_),
    .B(net4807),
    .Y(_01380_));
 NAND3x1_ASAP7_75t_R _07114_ (.A(_01376_),
    .B(_01379_),
    .C(net4807),
    .Y(_01381_));
 AOI22x1_ASAP7_75t_R _07115_ (.A1(_01372_),
    .A2(_01367_),
    .B1(_01380_),
    .B2(_01381_),
    .Y(_01382_));
 NAND3x1_ASAP7_75t_R _07116_ (.A(_01064_),
    .B(net4810),
    .C(_01042_),
    .Y(_01383_));
 INVx1_ASAP7_75t_R _07117_ (.A(_01042_),
    .Y(_01384_));
 INVx2_ASAP7_75t_R _07118_ (.A(_01064_),
    .Y(_01385_));
 INVx1_ASAP7_75t_R _07119_ (.A(net4810),
    .Y(_01386_));
 OAI21x1_ASAP7_75t_R _07120_ (.A1(_01384_),
    .A2(_01385_),
    .B(_01386_),
    .Y(_01387_));
 NOR2x1_ASAP7_75t_R _07121_ (.A(net5375),
    .B(net4808),
    .Y(_01388_));
 NAND2x1_ASAP7_75t_R _07122_ (.A(net4710),
    .B(_01388_),
    .Y(_01389_));
 NOR2x1_ASAP7_75t_R _07123_ (.A(net4649),
    .B(_01389_),
    .Y(_01390_));
 NAND2x1_ASAP7_75t_R _07124_ (.A(_01215_),
    .B(_01390_),
    .Y(_01391_));
 INVx1_ASAP7_75t_R _07125_ (.A(_01391_),
    .Y(_01392_));
 OAI21x1_ASAP7_75t_R _07126_ (.A1(net4583),
    .A2(net4591),
    .B(_01392_),
    .Y(_01393_));
 OAI21x1_ASAP7_75t_R _07127_ (.A1(net4811),
    .A2(net4833),
    .B(_00407_),
    .Y(_01394_));
 AOI21x1_ASAP7_75t_R _07128_ (.A1(net4708),
    .A2(net4709),
    .B(_01394_),
    .Y(_01395_));
 OAI21x1_ASAP7_75t_R _07129_ (.A1(net4645),
    .A2(net4648),
    .B(_01395_),
    .Y(_01396_));
 AOI21x1_ASAP7_75t_R _07130_ (.A1(_01390_),
    .A2(net4590),
    .B(_01396_),
    .Y(_01397_));
 NAND3x1_ASAP7_75t_R _07131_ (.A(_01393_),
    .B(net4812),
    .C(_01397_),
    .Y(_01398_));
 INVx1_ASAP7_75t_R _07132_ (.A(_01397_),
    .Y(_01399_));
 AOI21x1_ASAP7_75t_R _07133_ (.A1(net4536),
    .A2(net4535),
    .B(net4529),
    .Y(_01400_));
 INVx1_ASAP7_75t_R _07134_ (.A(net4812),
    .Y(_01401_));
 OAI21x1_ASAP7_75t_R _07135_ (.A1(_01399_),
    .A2(_01400_),
    .B(net4706),
    .Y(_01402_));
 AOI22x1_ASAP7_75t_R _07136_ (.A1(net4441),
    .A2(net4388),
    .B1(_01398_),
    .B2(_01402_),
    .Y(_01403_));
 NAND2x1_ASAP7_75t_R _07137_ (.A(_01382_),
    .B(_01403_),
    .Y(_01404_));
 NOR2x1_ASAP7_75t_R _07138_ (.A(_01404_),
    .B(_01357_),
    .Y(_01405_));
 NOR2x2_ASAP7_75t_R _07139_ (.A(_01286_),
    .B(_01283_),
    .Y(_01406_));
 NOR2x1_ASAP7_75t_R _07140_ (.A(_01305_),
    .B(_01302_),
    .Y(_01407_));
 NOR2x2_ASAP7_75t_R _07141_ (.A(_01406_),
    .B(_01407_),
    .Y(_01408_));
 INVx1_ASAP7_75t_R _07142_ (.A(_01300_),
    .Y(_01409_));
 INVx1_ASAP7_75t_R _07143_ (.A(_01297_),
    .Y(_01410_));
 NAND2x1_ASAP7_75t_R _07144_ (.A(_01409_),
    .B(_01410_),
    .Y(_01411_));
 OA21x2_ASAP7_75t_R _07145_ (.A1(_01253_),
    .A2(_01254_),
    .B(_01411_),
    .Y(_01412_));
 NAND2x1_ASAP7_75t_R _07146_ (.A(_01408_),
    .B(_01412_),
    .Y(_01413_));
 INVx2_ASAP7_75t_R _07147_ (.A(_01259_),
    .Y(_01414_));
 AOI21x1_ASAP7_75t_R _07148_ (.A1(_01274_),
    .A2(_01273_),
    .B(_01414_),
    .Y(_01415_));
 AOI22x1_ASAP7_75t_R _07149_ (.A1(_01228_),
    .A2(_01229_),
    .B1(_01279_),
    .B2(_01278_),
    .Y(_01416_));
 NAND2x1_ASAP7_75t_R _07150_ (.A(_01415_),
    .B(_01416_),
    .Y(_01417_));
 NOR2x1_ASAP7_75t_R _07151_ (.A(_01413_),
    .B(_01417_),
    .Y(_01418_));
 INVx1_ASAP7_75t_R _07152_ (.A(_01289_),
    .Y(_01419_));
 INVx1_ASAP7_75t_R _07153_ (.A(_01292_),
    .Y(_01420_));
 NOR2x1_ASAP7_75t_R _07154_ (.A(_01321_),
    .B(_01318_),
    .Y(_01421_));
 AOI21x1_ASAP7_75t_R _07155_ (.A1(_01419_),
    .A2(_01420_),
    .B(_01421_),
    .Y(_01422_));
 NAND2x1_ASAP7_75t_R _07156_ (.A(_01161_),
    .B(_01169_),
    .Y(_01423_));
 NAND2x1_ASAP7_75t_R _07157_ (.A(_01177_),
    .B(_01308_),
    .Y(_01424_));
 NOR2x1_ASAP7_75t_R _07158_ (.A(_01423_),
    .B(_01424_),
    .Y(_01425_));
 OA21x2_ASAP7_75t_R _07159_ (.A1(_01313_),
    .A2(_01316_),
    .B(_01309_),
    .Y(_01426_));
 NAND3x1_ASAP7_75t_R _07160_ (.A(_01422_),
    .B(_01425_),
    .C(_01426_),
    .Y(_01427_));
 NOR2x1_ASAP7_75t_R _07161_ (.A(_01427_),
    .B(_01157_),
    .Y(_01428_));
 NAND3x1_ASAP7_75t_R _07162_ (.A(_01428_),
    .B(_01405_),
    .C(_01418_),
    .Y(_01429_));
 NAND2x1_ASAP7_75t_R _07163_ (.A(_01067_),
    .B(_01012_),
    .Y(_01430_));
 NOR2x1_ASAP7_75t_R _07164_ (.A(net4647),
    .B(_01430_),
    .Y(_01431_));
 NAND2x1_ASAP7_75t_R _07165_ (.A(net4713),
    .B(_01039_),
    .Y(_01432_));
 AND2x2_ASAP7_75t_R _07166_ (.A(_01432_),
    .B(_01071_),
    .Y(_01433_));
 OAI21x1_ASAP7_75t_R _07167_ (.A1(net4646),
    .A2(_01430_),
    .B(_01433_),
    .Y(_01434_));
 AOI21x1_ASAP7_75t_R _07168_ (.A1(net4579),
    .A2(net4589),
    .B(_01434_),
    .Y(_01435_));
 NAND2x1_ASAP7_75t_R _07169_ (.A(_01232_),
    .B(_01431_),
    .Y(_01436_));
 AO21x1_ASAP7_75t_R _07170_ (.A1(_01285_),
    .A2(net5368),
    .B(_01436_),
    .Y(_01437_));
 AO21x1_ASAP7_75t_R _07171_ (.A1(_01435_),
    .A2(_01437_),
    .B(net4813),
    .Y(_01438_));
 NAND3x1_ASAP7_75t_R _07172_ (.A(_01435_),
    .B(net4813),
    .C(_01437_),
    .Y(_01439_));
 AND2x2_ASAP7_75t_R _07173_ (.A(_01438_),
    .B(_01439_),
    .Y(_01440_));
 INVx1_ASAP7_75t_R _07174_ (.A(net4383),
    .Y(_01441_));
 XOR2x2_ASAP7_75t_R _07175_ (.A(_01441_),
    .B(_01429_),
    .Y(_01442_));
 NOR2x1_ASAP7_75t_R _07176_ (.A(net4383),
    .B(net4286),
    .Y(_01443_));
 AOI21x1_ASAP7_75t_R _07177_ (.A1(_01442_),
    .A2(net4288),
    .B(_01443_),
    .Y(_01444_));
 OR5x1_ASAP7_75t_R _07178_ (.A(net4481),
    .B(_01293_),
    .C(_01322_),
    .D(_01327_),
    .E(_01324_),
    .Y(_01445_));
 NOR2x1_ASAP7_75t_R _07179_ (.A(_01306_),
    .B(_01260_),
    .Y(_01446_));
 AND3x1_ASAP7_75t_R _07180_ (.A(_01446_),
    .B(_01280_),
    .C(_01247_),
    .Y(_01447_));
 AOI22x1_ASAP7_75t_R _07181_ (.A1(_01340_),
    .A2(_01341_),
    .B1(_01211_),
    .B2(_01210_),
    .Y(_01448_));
 NAND2x1_ASAP7_75t_R _07182_ (.A(_01381_),
    .B(_01380_),
    .Y(_01449_));
 NAND2x1_ASAP7_75t_R _07183_ (.A(_01355_),
    .B(_01351_),
    .Y(_01450_));
 AND2x2_ASAP7_75t_R _07184_ (.A(_01450_),
    .B(_01449_),
    .Y(_01451_));
 NAND2x2_ASAP7_75t_R _07185_ (.A(_01448_),
    .B(_01451_),
    .Y(_01452_));
 NAND2x1p5_ASAP7_75t_R _07186_ (.A(_01383_),
    .B(_01387_),
    .Y(_01453_));
 NAND2x1_ASAP7_75t_R _07187_ (.A(_01367_),
    .B(_01372_),
    .Y(_01454_));
 AND2x4_ASAP7_75t_R _07188_ (.A(_01454_),
    .B(_01453_),
    .Y(_01455_));
 AOI22x1_ASAP7_75t_R _07189_ (.A1(_01439_),
    .A2(_01438_),
    .B1(_01402_),
    .B2(_01398_),
    .Y(_01456_));
 NAND2x1p5_ASAP7_75t_R _07190_ (.A(_01455_),
    .B(_01456_),
    .Y(_01457_));
 NOR2x1p5_ASAP7_75t_R _07191_ (.A(_01457_),
    .B(_01452_),
    .Y(_01458_));
 NAND2x1p5_ASAP7_75t_R _07192_ (.A(_01458_),
    .B(_01447_),
    .Y(_01459_));
 OAI21x1_ASAP7_75t_R _07193_ (.A1(_01459_),
    .A2(_01445_),
    .B(_01077_),
    .Y(_01460_));
 NAND2x1_ASAP7_75t_R _07194_ (.A(net4530),
    .B(_01362_),
    .Y(_01461_));
 AND3x1_ASAP7_75t_R _07195_ (.A(net4708),
    .B(_01068_),
    .C(_01401_),
    .Y(_01462_));
 INVx1_ASAP7_75t_R _07196_ (.A(net4834),
    .Y(_01463_));
 AOI21x1_ASAP7_75t_R _07197_ (.A1(_01401_),
    .A2(net4707),
    .B(_01463_),
    .Y(_01464_));
 OAI21x1_ASAP7_75t_R _07198_ (.A1(net4813),
    .A2(_01464_),
    .B(net4835),
    .Y(_01465_));
 AO21x1_ASAP7_75t_R _07199_ (.A1(_01461_),
    .A2(_01462_),
    .B(_01465_),
    .Y(_01466_));
 XOR2x2_ASAP7_75t_R _07200_ (.A(_01466_),
    .B(net4712),
    .Y(_01467_));
 XOR2x2_ASAP7_75t_R _07201_ (.A(net4333),
    .B(_01460_),
    .Y(_01468_));
 INVx3_ASAP7_75t_R _07202_ (.A(_01468_),
    .Y(_01469_));
 NAND2x1p5_ASAP7_75t_R _07203_ (.A(_01444_),
    .B(_01469_),
    .Y(_01470_));
 NAND2x1_ASAP7_75t_R _07204_ (.A(net4596),
    .B(net4597),
    .Y(_01471_));
 NOR2x1_ASAP7_75t_R _07205_ (.A(_01471_),
    .B(net4475),
    .Y(_01472_));
 INVx1_ASAP7_75t_R _07206_ (.A(net4474),
    .Y(_01473_));
 AND4x1_ASAP7_75t_R _07207_ (.A(_01426_),
    .B(net4598),
    .C(_01472_),
    .D(_01473_),
    .Y(_01474_));
 NAND2x1_ASAP7_75t_R _07208_ (.A(_01416_),
    .B(_01335_),
    .Y(_01475_));
 NAND2x1_ASAP7_75t_R _07209_ (.A(_01356_),
    .B(_01382_),
    .Y(_01476_));
 NOR2x1_ASAP7_75t_R _07210_ (.A(_01475_),
    .B(_01476_),
    .Y(_01477_));
 NAND2x1_ASAP7_75t_R _07211_ (.A(_01408_),
    .B(net5385),
    .Y(_01478_));
 NAND2x1_ASAP7_75t_R _07212_ (.A(_01415_),
    .B(_01412_),
    .Y(_01479_));
 NOR2x1_ASAP7_75t_R _07213_ (.A(_01478_),
    .B(_01479_),
    .Y(_01480_));
 AND2x2_ASAP7_75t_R _07214_ (.A(_01477_),
    .B(_01480_),
    .Y(_01481_));
 AOI21x1_ASAP7_75t_R _07215_ (.A1(_01474_),
    .A2(_01481_),
    .B(net4334),
    .Y(_01482_));
 INVx1_ASAP7_75t_R _07216_ (.A(net4334),
    .Y(_01483_));
 NAND3x1_ASAP7_75t_R _07217_ (.A(_01477_),
    .B(_01474_),
    .C(_01480_),
    .Y(_01484_));
 NOR2x1_ASAP7_75t_R _07218_ (.A(_01483_),
    .B(_01484_),
    .Y(_01485_));
 OAI21x1_ASAP7_75t_R _07219_ (.A1(_01482_),
    .A2(_01485_),
    .B(net4289),
    .Y(_01486_));
 NOR2x1_ASAP7_75t_R _07220_ (.A(_01483_),
    .B(net4286),
    .Y(_01487_));
 INVx1_ASAP7_75t_R _07221_ (.A(_01487_),
    .Y(_01488_));
 INVx1_ASAP7_75t_R _07222_ (.A(net4481),
    .Y(_01489_));
 NAND2x1_ASAP7_75t_R _07223_ (.A(_01489_),
    .B(net4443),
    .Y(_01490_));
 INVx1_ASAP7_75t_R _07224_ (.A(_01490_),
    .Y(_01491_));
 NOR2x1_ASAP7_75t_R _07225_ (.A(net4444),
    .B(_01293_),
    .Y(_01492_));
 NAND2x1_ASAP7_75t_R _07226_ (.A(_01492_),
    .B(_01446_),
    .Y(_01493_));
 NAND2x1_ASAP7_75t_R _07227_ (.A(_01280_),
    .B(_01247_),
    .Y(_01494_));
 NOR3x1_ASAP7_75t_R _07228_ (.A(net4234),
    .B(_01493_),
    .C(_01494_),
    .Y(_01495_));
 AOI21x1_ASAP7_75t_R _07229_ (.A1(_01491_),
    .A2(_01495_),
    .B(net4340),
    .Y(_01496_));
 INVx1_ASAP7_75t_R _07230_ (.A(net4380),
    .Y(_01497_));
 XOR2x2_ASAP7_75t_R _07231_ (.A(_01496_),
    .B(_01497_),
    .Y(_01498_));
 AND2x2_ASAP7_75t_R _07232_ (.A(_01455_),
    .B(_01451_),
    .Y(_01499_));
 NAND2x1_ASAP7_75t_R _07233_ (.A(_01247_),
    .B(net4433),
    .Y(_01500_));
 NOR3x1_ASAP7_75t_R _07234_ (.A(_01281_),
    .B(_01329_),
    .C(_01500_),
    .Y(_01501_));
 AOI21x1_ASAP7_75t_R _07235_ (.A1(_01499_),
    .A2(_01501_),
    .B(net4340),
    .Y(_01502_));
 AND2x2_ASAP7_75t_R _07236_ (.A(_01398_),
    .B(_01402_),
    .Y(_01503_));
 XOR2x2_ASAP7_75t_R _07237_ (.A(_01502_),
    .B(_01503_),
    .Y(_01504_));
 AOI211x1_ASAP7_75t_R _07238_ (.A1(_01486_),
    .A2(_01488_),
    .B(_01498_),
    .C(_01504_),
    .Y(_01505_));
 INVx1_ASAP7_75t_R _07239_ (.A(_01403_),
    .Y(_01506_));
 OR3x1_ASAP7_75t_R _07240_ (.A(_01467_),
    .B(_01440_),
    .C(_01506_),
    .Y(_01507_));
 NOR2x1_ASAP7_75t_R _07241_ (.A(_01476_),
    .B(_01507_),
    .Y(_01508_));
 AND5x1_ASAP7_75t_R _07242_ (.A(net4434),
    .B(_01170_),
    .C(net5385),
    .D(_01408_),
    .E(_01473_),
    .Y(_01509_));
 NOR2x1_ASAP7_75t_R _07243_ (.A(net4283),
    .B(net4379),
    .Y(_01510_));
 AND4x1_ASAP7_75t_R _07244_ (.A(_01508_),
    .B(net4286),
    .C(_01509_),
    .D(_01510_),
    .Y(_01511_));
 NAND2x1p5_ASAP7_75t_R _07245_ (.A(_01468_),
    .B(_01511_),
    .Y(_01512_));
 OAI21x1_ASAP7_75t_R _07246_ (.A1(_01470_),
    .A2(_01505_),
    .B(_01512_),
    .Y(_01513_));
 INVx1_ASAP7_75t_R _07247_ (.A(net4054),
    .Y(_01514_));
 XOR2x2_ASAP7_75t_R _07248_ (.A(_01513_),
    .B(_01514_),
    .Y(_01515_));
 INVx1_ASAP7_75t_R _07249_ (.A(net3975),
    .Y(_01516_));
 NAND2x1_ASAP7_75t_R _07250_ (.A(net4175),
    .B(net4055),
    .Y(_01517_));
 NAND2x1_ASAP7_75t_R _07251_ (.A(_01469_),
    .B(_01511_),
    .Y(_01518_));
 NAND2x1_ASAP7_75t_R _07252_ (.A(_01517_),
    .B(_01518_),
    .Y(_01519_));
 INVx2_ASAP7_75t_R _07253_ (.A(_01519_),
    .Y(_01520_));
 NAND2x1_ASAP7_75t_R _07254_ (.A(net3974),
    .B(_01515_),
    .Y(_01521_));
 XOR2x2_ASAP7_75t_R _07255_ (.A(_01429_),
    .B(net4383),
    .Y(_01522_));
 INVx1_ASAP7_75t_R _07256_ (.A(_01443_),
    .Y(_01523_));
 OAI21x1_ASAP7_75t_R _07257_ (.A1(net4341),
    .A2(_01522_),
    .B(_01523_),
    .Y(_01524_));
 XNOR2x2_ASAP7_75t_R _07258_ (.A(_01503_),
    .B(_01502_),
    .Y(_01525_));
 AO21x1_ASAP7_75t_R _07259_ (.A1(_01511_),
    .A2(_01469_),
    .B(_01525_),
    .Y(_01526_));
 OR3x1_ASAP7_75t_R _07260_ (.A(_01513_),
    .B(net4053),
    .C(_01526_),
    .Y(_01527_));
 INVx1_ASAP7_75t_R _07261_ (.A(_01527_),
    .Y(_01528_));
 INVx1_ASAP7_75t_R _07262_ (.A(_01486_),
    .Y(_01529_));
 OAI21x1_ASAP7_75t_R _07263_ (.A1(net4233),
    .A2(_01529_),
    .B(_01525_),
    .Y(_01530_));
 NOR2x1_ASAP7_75t_R _07264_ (.A(_01468_),
    .B(_01524_),
    .Y(_01531_));
 OAI21x1_ASAP7_75t_R _07265_ (.A1(net4054),
    .A2(_01530_),
    .B(_01531_),
    .Y(_01532_));
 OR2x2_ASAP7_75t_R _07266_ (.A(_01444_),
    .B(_01530_),
    .Y(_01533_));
 INVx1_ASAP7_75t_R _07267_ (.A(net4434),
    .Y(_01534_));
 INVx1_ASAP7_75t_R _07268_ (.A(net4534),
    .Y(_01535_));
 INVx1_ASAP7_75t_R _07269_ (.A(net4537),
    .Y(_01536_));
 OR3x1_ASAP7_75t_R _07270_ (.A(_01171_),
    .B(_01535_),
    .C(_01536_),
    .Y(_01537_));
 NOR2x1_ASAP7_75t_R _07271_ (.A(net4377),
    .B(_01537_),
    .Y(_01538_));
 NAND3x1_ASAP7_75t_R _07272_ (.A(_01538_),
    .B(net4384),
    .C(net4387),
    .Y(_01539_));
 INVx1_ASAP7_75t_R _07273_ (.A(net4438),
    .Y(_01540_));
 NOR3x1_ASAP7_75t_R _07274_ (.A(_01539_),
    .B(_01540_),
    .C(net4283),
    .Y(_01541_));
 INVx1_ASAP7_75t_R _07275_ (.A(net4284),
    .Y(_01542_));
 NAND3x1_ASAP7_75t_R _07276_ (.A(_01541_),
    .B(net4231),
    .C(net4389),
    .Y(_01543_));
 AND3x1_ASAP7_75t_R _07277_ (.A(_01077_),
    .B(_01441_),
    .C(_01403_),
    .Y(_01544_));
 INVx1_ASAP7_75t_R _07278_ (.A(_01544_),
    .Y(_01545_));
 NOR3x1_ASAP7_75t_R _07279_ (.A(_01543_),
    .B(net4333),
    .C(_01545_),
    .Y(_01546_));
 AOI21x1_ASAP7_75t_R _07280_ (.A1(_01533_),
    .A2(_01546_),
    .B(net4026),
    .Y(_01547_));
 NAND2x2_ASAP7_75t_R _07281_ (.A(net3991),
    .B(_01547_),
    .Y(_01548_));
 INVx2_ASAP7_75t_R _07282_ (.A(_01548_),
    .Y(_01549_));
 AND5x1_ASAP7_75t_R _07283_ (.A(net4761),
    .B(net4435),
    .C(net4596),
    .D(_01145_),
    .E(net4597),
    .Y(_01550_));
 AND4x1_ASAP7_75t_R _07284_ (.A(net4337),
    .B(net4434),
    .C(net5385),
    .D(net4387),
    .Y(_01551_));
 INVx1_ASAP7_75t_R _07285_ (.A(net4336),
    .Y(_01552_));
 AND5x1_ASAP7_75t_R _07286_ (.A(_01550_),
    .B(net5143),
    .C(_01551_),
    .D(_01542_),
    .E(_01552_),
    .Y(_01553_));
 INVx1_ASAP7_75t_R _07287_ (.A(net4381),
    .Y(_01554_));
 XOR2x2_ASAP7_75t_R _07288_ (.A(_01553_),
    .B(_01554_),
    .Y(_01555_));
 NOR2x1_ASAP7_75t_R _07289_ (.A(net4332),
    .B(net4290),
    .Y(_01556_));
 AO21x1_ASAP7_75t_R _07290_ (.A1(_01555_),
    .A2(net4290),
    .B(_01556_),
    .Y(_01557_));
 BUFx3_ASAP7_75t_R place3023 (.A(_03954_),
    .Y(net3023));
 INVx1_ASAP7_75t_R _07292_ (.A(net4051),
    .Y(_01559_));
 AOI211x1_ASAP7_75t_R _07293_ (.A1(_01521_),
    .A2(_01528_),
    .B(_01549_),
    .C(_01559_),
    .Y(_01560_));
 OAI21x1_ASAP7_75t_R _07294_ (.A1(_01559_),
    .A2(_01521_),
    .B(_01528_),
    .Y(_01561_));
 AOI21x1_ASAP7_75t_R _07295_ (.A1(net3971),
    .A2(_01561_),
    .B(net4052),
    .Y(_01562_));
 NOR2x1_ASAP7_75t_R _07296_ (.A(net4341),
    .B(net4282),
    .Y(_01563_));
 XOR2x2_ASAP7_75t_R _07297_ (.A(_01563_),
    .B(net4335),
    .Y(_01564_));
 OAI21x1_ASAP7_75t_R _07298_ (.A1(_01562_),
    .A2(_01560_),
    .B(_01564_),
    .Y(_01565_));
 NOR2x2_ASAP7_75t_R _07299_ (.A(_01516_),
    .B(_01565_),
    .Y(_01566_));
 NOR2x1_ASAP7_75t_R _07300_ (.A(_01514_),
    .B(_01513_),
    .Y(_01567_));
 AOI21x1_ASAP7_75t_R _07301_ (.A1(net4001),
    .A2(_01532_),
    .B(net4054),
    .Y(_01568_));
 NOR3x1_ASAP7_75t_R _07302_ (.A(_01567_),
    .B(_01568_),
    .C(net3985),
    .Y(_01569_));
 AOI22x1_ASAP7_75t_R _07303_ (.A1(_01569_),
    .A2(net4051),
    .B1(_01548_),
    .B2(net3972),
    .Y(_01570_));
 INVx1_ASAP7_75t_R _07304_ (.A(_01526_),
    .Y(_01571_));
 NAND2x1_ASAP7_75t_R _07305_ (.A(net3973),
    .B(_01568_),
    .Y(_01572_));
 INVx1_ASAP7_75t_R _07306_ (.A(net4337),
    .Y(_01573_));
 INVx1_ASAP7_75t_R _07307_ (.A(net4384),
    .Y(_01574_));
 OR4x1_ASAP7_75t_R _07308_ (.A(_01171_),
    .B(_01535_),
    .C(_01536_),
    .D(_01534_),
    .Y(_01575_));
 NOR2x1_ASAP7_75t_R _07309_ (.A(_01574_),
    .B(_01575_),
    .Y(_01576_));
 NAND2x1_ASAP7_75t_R _07310_ (.A(net4387),
    .B(_01576_),
    .Y(_01577_));
 NOR2x1_ASAP7_75t_R _07311_ (.A(_01573_),
    .B(_01577_),
    .Y(_01578_));
 AND3x1_ASAP7_75t_R _07312_ (.A(net4389),
    .B(_01335_),
    .C(_01356_),
    .Y(_01579_));
 AND4x1_ASAP7_75t_R _07313_ (.A(_01578_),
    .B(net4438),
    .C(net4385),
    .D(_01579_),
    .Y(_01580_));
 NAND2x1_ASAP7_75t_R _07314_ (.A(net4230),
    .B(_01580_),
    .Y(_01581_));
 AOI211x1_ASAP7_75t_R _07315_ (.A1(net3990),
    .A2(net4002),
    .B(_01581_),
    .C(net4333),
    .Y(_01582_));
 AO21x1_ASAP7_75t_R _07316_ (.A1(_01571_),
    .A2(_01572_),
    .B(_01582_),
    .Y(_01583_));
 XOR2x2_ASAP7_75t_R _07317_ (.A(_01570_),
    .B(_01583_),
    .Y(_01584_));
 AOI21x1_ASAP7_75t_R _07318_ (.A1(net4051),
    .A2(_01569_),
    .B(net3972),
    .Y(_01585_));
 XOR2x2_ASAP7_75t_R _07319_ (.A(_01568_),
    .B(net3985),
    .Y(_01586_));
 NOR3x1_ASAP7_75t_R _07320_ (.A(_01585_),
    .B(net3964),
    .C(_01586_),
    .Y(_01587_));
 NAND2x2_ASAP7_75t_R _07321_ (.A(_01515_),
    .B(net4051),
    .Y(_01588_));
 XOR2x2_ASAP7_75t_R _07322_ (.A(_01568_),
    .B(_01520_),
    .Y(_01589_));
 XOR2x1_ASAP7_75t_R _07323_ (.A(_01588_),
    .Y(_01590_),
    .B(_01589_));
 NAND3x1_ASAP7_75t_R _07324_ (.A(_01515_),
    .B(net4051),
    .C(net3974),
    .Y(_01591_));
 AOI21x1_ASAP7_75t_R _07325_ (.A1(_01528_),
    .A2(_01591_),
    .B(_01549_),
    .Y(_01592_));
 NOR2x1_ASAP7_75t_R _07326_ (.A(_01592_),
    .B(_01590_),
    .Y(_01593_));
 NOR2x1_ASAP7_75t_R _07327_ (.A(_01587_),
    .B(_01593_),
    .Y(_01594_));
 NAND2x1_ASAP7_75t_R _07328_ (.A(_01594_),
    .B(_01584_),
    .Y(_01595_));
 NAND2x1_ASAP7_75t_R _07329_ (.A(_01583_),
    .B(_01570_),
    .Y(_01596_));
 NAND2x1_ASAP7_75t_R _07330_ (.A(net4056),
    .B(net3991),
    .Y(_01597_));
 AO21x1_ASAP7_75t_R _07331_ (.A1(_01596_),
    .A2(_01597_),
    .B(net3953),
    .Y(_01598_));
 OAI21x1_ASAP7_75t_R _07332_ (.A1(_01566_),
    .A2(_01595_),
    .B(_01598_),
    .Y(_01599_));
 INVx1_ASAP7_75t_R _07333_ (.A(_01564_),
    .Y(_01600_));
 OAI21x1_ASAP7_75t_R _07334_ (.A1(net3965),
    .A2(net3953),
    .B(net4025),
    .Y(_01601_));
 INVx1_ASAP7_75t_R _07335_ (.A(_01560_),
    .Y(_01602_));
 NAND2x1_ASAP7_75t_R _07336_ (.A(_01601_),
    .B(_01602_),
    .Y(_01603_));
 NOR2x1_ASAP7_75t_R _07337_ (.A(net4100),
    .B(_01603_),
    .Y(_01604_));
 INVx1_ASAP7_75t_R _07338_ (.A(_01603_),
    .Y(_01605_));
 NOR2x1_ASAP7_75t_R _07339_ (.A(net4174),
    .B(_01605_),
    .Y(_01606_));
 OR2x2_ASAP7_75t_R _07340_ (.A(_01604_),
    .B(_01606_),
    .Y(_01607_));
 NOR2x1_ASAP7_75t_R _07341_ (.A(net3926),
    .B(_01599_),
    .Y(_01608_));
 AO21x1_ASAP7_75t_R _07342_ (.A1(_01599_),
    .A2(_01607_),
    .B(_01608_),
    .Y(_01609_));
 AOI21x1_ASAP7_75t_R _07343_ (.A1(_01598_),
    .A2(_01595_),
    .B(net3927),
    .Y(_01610_));
 XOR2x2_ASAP7_75t_R _07344_ (.A(_01610_),
    .B(net3936),
    .Y(_01611_));
 INVx1_ASAP7_75t_R _07345_ (.A(net3952),
    .Y(_01612_));
 XOR2x2_ASAP7_75t_R _07346_ (.A(net3975),
    .B(_01559_),
    .Y(_01613_));
 AO21x1_ASAP7_75t_R _07347_ (.A1(_01561_),
    .A2(net3971),
    .B(_01613_),
    .Y(_01614_));
 OAI21x1_ASAP7_75t_R _07348_ (.A1(_01516_),
    .A2(_01612_),
    .B(_01614_),
    .Y(_01615_));
 INVx1_ASAP7_75t_R _07349_ (.A(net3934),
    .Y(_01616_));
 NOR2x1p5_ASAP7_75t_R _07350_ (.A(_01599_),
    .B(_01616_),
    .Y(_01617_));
 XOR2x2_ASAP7_75t_R _07351_ (.A(_01615_),
    .B(_01565_),
    .Y(_01618_));
 AOI21x1_ASAP7_75t_R _07352_ (.A1(_01601_),
    .A2(_01602_),
    .B(_01600_),
    .Y(_01619_));
 NAND2x1_ASAP7_75t_R _07353_ (.A(net3975),
    .B(_01619_),
    .Y(_01620_));
 INVx1_ASAP7_75t_R _07354_ (.A(_01584_),
    .Y(_01621_));
 NAND2x1_ASAP7_75t_R _07355_ (.A(net3963),
    .B(net3952),
    .Y(_01622_));
 XOR2x2_ASAP7_75t_R _07356_ (.A(_01588_),
    .B(_01586_),
    .Y(_01623_));
 OAI21x1_ASAP7_75t_R _07357_ (.A1(net3965),
    .A2(net3953),
    .B(_01623_),
    .Y(_01624_));
 NAND2x1_ASAP7_75t_R _07358_ (.A(_01622_),
    .B(_01624_),
    .Y(_01625_));
 NOR2x1_ASAP7_75t_R _07359_ (.A(_01621_),
    .B(_01625_),
    .Y(_01626_));
 INVx1_ASAP7_75t_R _07360_ (.A(_01598_),
    .Y(_01627_));
 AOI21x1_ASAP7_75t_R _07361_ (.A1(_01620_),
    .A2(_01626_),
    .B(_01627_),
    .Y(_01628_));
 NOR2x1_ASAP7_75t_R _07362_ (.A(_01618_),
    .B(_01628_),
    .Y(_01629_));
 NOR2x2_ASAP7_75t_R _07363_ (.A(_01629_),
    .B(_01617_),
    .Y(_01630_));
 NAND2x2_ASAP7_75t_R _07364_ (.A(_01611_),
    .B(_01630_),
    .Y(_01631_));
 NOR2x1_ASAP7_75t_R _07365_ (.A(_01625_),
    .B(net3927),
    .Y(_01632_));
 AO21x1_ASAP7_75t_R _07366_ (.A1(_01632_),
    .A2(_01627_),
    .B(_01584_),
    .Y(_01633_));
 NAND2x1_ASAP7_75t_R _07367_ (.A(net3923),
    .B(net3922),
    .Y(_01634_));
 AND2x2_ASAP7_75t_R _07368_ (.A(_01633_),
    .B(_01634_),
    .Y(_01635_));
 INVx1_ASAP7_75t_R _07369_ (.A(_01635_),
    .Y(_01636_));
 OAI21x1_ASAP7_75t_R _07370_ (.A1(_01609_),
    .A2(_01631_),
    .B(_01636_),
    .Y(_01637_));
 NAND2x1_ASAP7_75t_R _07371_ (.A(net4477),
    .B(net4478),
    .Y(_01638_));
 INVx1_ASAP7_75t_R _07372_ (.A(net4442),
    .Y(_01639_));
 NOR2x1_ASAP7_75t_R _07373_ (.A(net4341),
    .B(net4232),
    .Y(_01640_));
 AO21x1_ASAP7_75t_R _07374_ (.A1(net4288),
    .A2(_01639_),
    .B(_01640_),
    .Y(_01641_));
 XNOR2x2_ASAP7_75t_R _07375_ (.A(_01638_),
    .B(_01641_),
    .Y(_01642_));
 XOR2x2_ASAP7_75t_R _07376_ (.A(net4100),
    .B(_01599_),
    .Y(_01643_));
 NOR2x2_ASAP7_75t_R _07377_ (.A(net4050),
    .B(_01643_),
    .Y(_01644_));
 NAND3x1_ASAP7_75t_R _07378_ (.A(_01637_),
    .B(net3894),
    .C(_01644_),
    .Y(_01645_));
 INVx1_ASAP7_75t_R _07379_ (.A(_01644_),
    .Y(_01646_));
 INVx1_ASAP7_75t_R _07380_ (.A(_01637_),
    .Y(_01647_));
 INVx1_ASAP7_75t_R _07381_ (.A(net3894),
    .Y(_01648_));
 OAI21x1_ASAP7_75t_R _07382_ (.A1(_01646_),
    .A2(_01647_),
    .B(_01648_),
    .Y(_01649_));
 NAND2x1_ASAP7_75t_R _07383_ (.A(net3934),
    .B(net3915),
    .Y(_01650_));
 OAI21x1_ASAP7_75t_R _07384_ (.A1(net3915),
    .A2(net3924),
    .B(_01650_),
    .Y(_01651_));
 AOI22x1_ASAP7_75t_R _07385_ (.A1(_01631_),
    .A2(_01636_),
    .B1(_01644_),
    .B2(net3935),
    .Y(_01652_));
 NAND2x1_ASAP7_75t_R _07386_ (.A(_01651_),
    .B(_01652_),
    .Y(_01653_));
 INVx3_ASAP7_75t_R _07387_ (.A(_01631_),
    .Y(_01654_));
 XOR2x2_ASAP7_75t_R _07388_ (.A(net4174),
    .B(_01599_),
    .Y(_01655_));
 INVx1_ASAP7_75t_R _07389_ (.A(_01642_),
    .Y(_01656_));
 NAND3x2_ASAP7_75t_R _07390_ (.B(_01655_),
    .C(net3935),
    .Y(_01657_),
    .A(_01656_));
 OAI21x1_ASAP7_75t_R _07391_ (.A1(net3892),
    .A2(_01654_),
    .B(_01657_),
    .Y(_01658_));
 NAND2x1_ASAP7_75t_R _07392_ (.A(net3893),
    .B(_01658_),
    .Y(_01659_));
 AOI22x1_ASAP7_75t_R _07393_ (.A1(_01645_),
    .A2(_01649_),
    .B1(_01653_),
    .B2(_01659_),
    .Y(_01660_));
 AND2x2_ASAP7_75t_R _07394_ (.A(_01607_),
    .B(_01599_),
    .Y(_01661_));
 OAI21x1_ASAP7_75t_R _07395_ (.A1(_01608_),
    .A2(_01661_),
    .B(net3925),
    .Y(_01662_));
 OAI21x1_ASAP7_75t_R _07396_ (.A1(net4050),
    .A2(_01643_),
    .B(_01611_),
    .Y(_01663_));
 NOR2x1_ASAP7_75t_R _07397_ (.A(_01662_),
    .B(_01663_),
    .Y(_01664_));
 OAI21x1_ASAP7_75t_R _07398_ (.A1(_01664_),
    .A2(_01637_),
    .B(net4050),
    .Y(_01665_));
 AOI21x1_ASAP7_75t_R _07399_ (.A1(_01657_),
    .A2(_01654_),
    .B(net3892),
    .Y(_01666_));
 NAND2x2_ASAP7_75t_R _07400_ (.A(_01666_),
    .B(net4024),
    .Y(_01667_));
 AOI21x1_ASAP7_75t_R _07401_ (.A1(_01665_),
    .A2(_01667_),
    .B(_01333_),
    .Y(_01668_));
 NAND2x1p5_ASAP7_75t_R _07402_ (.A(net3905),
    .B(_01668_),
    .Y(_01669_));
 NAND2x1_ASAP7_75t_R _07403_ (.A(net3893),
    .B(_01657_),
    .Y(_01670_));
 INVx1_ASAP7_75t_R _07404_ (.A(_01611_),
    .Y(_01671_));
 OA21x2_ASAP7_75t_R _07405_ (.A1(_01670_),
    .A2(_01636_),
    .B(_01671_),
    .Y(_01672_));
 AOI21x1_ASAP7_75t_R _07406_ (.A1(net3891),
    .A2(net3871),
    .B(_01672_),
    .Y(_01673_));
 AOI21x1_ASAP7_75t_R _07407_ (.A1(_01660_),
    .A2(_01669_),
    .B(net5399),
    .Y(_01674_));
 NAND2x1p5_ASAP7_75t_R _07408_ (.A(net4101),
    .B(_01674_),
    .Y(_01675_));
 NAND2x1_ASAP7_75t_R _07409_ (.A(_01659_),
    .B(_01653_),
    .Y(_01676_));
 NAND2x1_ASAP7_75t_R _07410_ (.A(_01649_),
    .B(_01645_),
    .Y(_01677_));
 NAND2x1_ASAP7_75t_R _07411_ (.A(_01676_),
    .B(_01677_),
    .Y(_01678_));
 AOI211x1_ASAP7_75t_R _07412_ (.A1(_01667_),
    .A2(_01665_),
    .B(net3906),
    .C(net4176),
    .Y(_01679_));
 INVx1_ASAP7_75t_R _07413_ (.A(_01673_),
    .Y(_01680_));
 OAI21x1_ASAP7_75t_R _07414_ (.A1(_01679_),
    .A2(_01678_),
    .B(_01680_),
    .Y(_01681_));
 NAND2x1_ASAP7_75t_R _07415_ (.A(net4176),
    .B(_01681_),
    .Y(_01682_));
 NAND2x1_ASAP7_75t_R _07416_ (.A(net3795),
    .B(net3794),
    .Y(_01683_));
 INVx1_ASAP7_75t_R _07417_ (.A(_01683_),
    .Y(_01684_));
 NAND2x1_ASAP7_75t_R _07418_ (.A(net4488),
    .B(net4489),
    .Y(_01685_));
 XNOR2x2_ASAP7_75t_R _07419_ (.A(_01685_),
    .B(net4173),
    .Y(_01686_));
 OAI21x1_ASAP7_75t_R _07420_ (.A1(net3860),
    .A2(_01660_),
    .B(_01669_),
    .Y(_01687_));
 XOR2x2_ASAP7_75t_R _07421_ (.A(net5888),
    .B(net3831),
    .Y(_01688_));
 OAI21x1_ASAP7_75t_R _07422_ (.A1(net4050),
    .A2(net3861),
    .B(net3906),
    .Y(_01689_));
 OA21x2_ASAP7_75t_R _07423_ (.A1(_01646_),
    .A2(net3861),
    .B(_01689_),
    .Y(_01690_));
 XNOR2x2_ASAP7_75t_R _07424_ (.A(net3833),
    .B(_01690_),
    .Y(_01691_));
 NAND2x1_ASAP7_75t_R _07425_ (.A(_01674_),
    .B(net3830),
    .Y(_01692_));
 OAI21x1_ASAP7_75t_R _07426_ (.A1(_01691_),
    .A2(net5766),
    .B(_01692_),
    .Y(_01693_));
 NOR2x1p5_ASAP7_75t_R _07427_ (.A(_01688_),
    .B(_01693_),
    .Y(_01694_));
 INVx1_ASAP7_75t_R _07428_ (.A(_01686_),
    .Y(_01695_));
 NAND2x1_ASAP7_75t_R _07429_ (.A(net3862),
    .B(net3849),
    .Y(_01696_));
 INVx1_ASAP7_75t_R _07430_ (.A(net3829),
    .Y(_01697_));
 AOI21x1_ASAP7_75t_R _07431_ (.A1(_01675_),
    .A2(_01682_),
    .B(_01697_),
    .Y(_01698_));
 NAND2x1p5_ASAP7_75t_R _07432_ (.A(_01695_),
    .B(_01698_),
    .Y(_01699_));
 INVx1_ASAP7_75t_R _07433_ (.A(_01676_),
    .Y(_01700_));
 INVx1_ASAP7_75t_R _07434_ (.A(_01677_),
    .Y(_01701_));
 AOI211x1_ASAP7_75t_R _07435_ (.A1(_01680_),
    .A2(_01700_),
    .B(net5455),
    .C(_01701_),
    .Y(_01702_));
 XOR2x2_ASAP7_75t_R _07436_ (.A(_01702_),
    .B(net3832),
    .Y(_01703_));
 AOI21x1_ASAP7_75t_R _07437_ (.A1(_01694_),
    .A2(_01699_),
    .B(_01703_),
    .Y(_01704_));
 NAND2x2_ASAP7_75t_R _07438_ (.A(_01704_),
    .B(net4099),
    .Y(_01705_));
 NOR2x1_ASAP7_75t_R _07439_ (.A(net4341),
    .B(net4285),
    .Y(_01706_));
 NAND2x1_ASAP7_75t_R _07440_ (.A(net4490),
    .B(net4491),
    .Y(_01707_));
 INVx1_ASAP7_75t_R _07441_ (.A(_01707_),
    .Y(_01708_));
 XOR2x2_ASAP7_75t_R _07442_ (.A(_01706_),
    .B(_01708_),
    .Y(_01709_));
 INVx1_ASAP7_75t_R _07443_ (.A(_01709_),
    .Y(_01710_));
 AND3x1_ASAP7_75t_R _07444_ (.A(net5400),
    .B(net3905),
    .C(net3833),
    .Y(_01711_));
 AOI21x1_ASAP7_75t_R _07445_ (.A1(net3833),
    .A2(net3805),
    .B(net3830),
    .Y(_01712_));
 XOR2x2_ASAP7_75t_R _07446_ (.A(_01701_),
    .B(_01687_),
    .Y(_01713_));
 OAI21x1_ASAP7_75t_R _07447_ (.A1(_01711_),
    .A2(_01712_),
    .B(_01713_),
    .Y(_01714_));
 NOR2x1_ASAP7_75t_R _07448_ (.A(_01698_),
    .B(_01714_),
    .Y(_01715_));
 OAI21x1_ASAP7_75t_R _07449_ (.A1(net3793),
    .A2(_01715_),
    .B(net4049),
    .Y(_01716_));
 NAND3x2_ASAP7_75t_R _07450_ (.B(_01705_),
    .C(_01710_),
    .Y(_01717_),
    .A(_01716_));
 XOR2x2_ASAP7_75t_R _07451_ (.A(_01696_),
    .B(_01334_),
    .Y(_01718_));
 NAND2x1_ASAP7_75t_R _07452_ (.A(_01718_),
    .B(net3805),
    .Y(_01719_));
 OAI21x1_ASAP7_75t_R _07453_ (.A1(_01697_),
    .A2(net5889),
    .B(_01719_),
    .Y(_01720_));
 INVx1_ASAP7_75t_R _07454_ (.A(net3772),
    .Y(_01721_));
 NAND2x1p5_ASAP7_75t_R _07455_ (.A(_01721_),
    .B(_01704_),
    .Y(_01722_));
 AO21x1_ASAP7_75t_R _07456_ (.A1(net5437),
    .A2(net3862),
    .B(net3906),
    .Y(_01723_));
 AOI211x1_ASAP7_75t_R _07457_ (.A1(_01660_),
    .A2(_01723_),
    .B(net5400),
    .C(net4176),
    .Y(_01724_));
 NOR2x1p5_ASAP7_75t_R _07458_ (.A(net4101),
    .B(_01674_),
    .Y(_01725_));
 OAI21x1_ASAP7_75t_R _07459_ (.A1(net3818),
    .A2(_01725_),
    .B(_01695_),
    .Y(_01726_));
 XOR2x2_ASAP7_75t_R _07460_ (.A(_01726_),
    .B(_01720_),
    .Y(_01727_));
 OAI21x1_ASAP7_75t_R _07461_ (.A1(_01724_),
    .A2(_01725_),
    .B(net3829),
    .Y(_01728_));
 NOR2x1_ASAP7_75t_R _07462_ (.A(net4099),
    .B(_01728_),
    .Y(_01729_));
 INVx1_ASAP7_75t_R _07463_ (.A(_01703_),
    .Y(_01730_));
 OAI21x1_ASAP7_75t_R _07464_ (.A1(_01714_),
    .A2(_01729_),
    .B(_01730_),
    .Y(_01731_));
 NAND2x1_ASAP7_75t_R _07465_ (.A(_01727_),
    .B(_01731_),
    .Y(_01732_));
 AOI21x1_ASAP7_75t_R _07466_ (.A1(net3773),
    .A2(_01730_),
    .B(_01729_),
    .Y(_01733_));
 NAND2x1_ASAP7_75t_R _07467_ (.A(net3774),
    .B(_01733_),
    .Y(_01734_));
 INVx1_ASAP7_75t_R _07468_ (.A(net3774),
    .Y(_01735_));
 OAI21x1_ASAP7_75t_R _07469_ (.A1(net3792),
    .A2(_01694_),
    .B(_01699_),
    .Y(_01736_));
 NAND2x1_ASAP7_75t_R _07470_ (.A(_01735_),
    .B(_01736_),
    .Y(_01737_));
 AOI22x1_ASAP7_75t_R _07471_ (.A1(_01732_),
    .A2(_01722_),
    .B1(_01734_),
    .B2(_01737_),
    .Y(_01738_));
 OAI21x1_ASAP7_75t_R _07472_ (.A1(_01717_),
    .A2(net3761),
    .B(_01738_),
    .Y(_01739_));
 NOR2x1_ASAP7_75t_R _07473_ (.A(net3774),
    .B(_01729_),
    .Y(_01740_));
 AO21x1_ASAP7_75t_R _07474_ (.A1(_01740_),
    .A2(_01703_),
    .B(net5438),
    .Y(_01741_));
 NAND2x1_ASAP7_75t_R _07475_ (.A(_01694_),
    .B(net3760),
    .Y(_01742_));
 AND2x2_ASAP7_75t_R _07476_ (.A(_01741_),
    .B(_01742_),
    .Y(_01743_));
 INVx2_ASAP7_75t_R _07477_ (.A(_01743_),
    .Y(_01744_));
 NAND2x1_ASAP7_75t_R _07478_ (.A(net3745),
    .B(_01722_),
    .Y(_01745_));
 OAI21x1_ASAP7_75t_R _07479_ (.A1(net3761),
    .A2(net3730),
    .B(net3725),
    .Y(_01746_));
 NAND2x1_ASAP7_75t_R _07480_ (.A(net3743),
    .B(net3744),
    .Y(_01747_));
 INVx1_ASAP7_75t_R _07481_ (.A(net3724),
    .Y(_01748_));
 OAI21x1_ASAP7_75t_R _07482_ (.A1(_01744_),
    .A2(_01746_),
    .B(_01748_),
    .Y(_01749_));
 NAND2x2_ASAP7_75t_R _07483_ (.A(net3715),
    .B(_01749_),
    .Y(_01750_));
 INVx2_ASAP7_75t_R _07484_ (.A(_01750_),
    .Y(_01751_));
 NAND3x1_ASAP7_75t_R _07485_ (.A(net5763),
    .B(net3775),
    .C(_01716_),
    .Y(_01752_));
 AOI211x1_ASAP7_75t_R _07486_ (.A1(_01738_),
    .A2(_01752_),
    .B(_01743_),
    .C(net4172),
    .Y(_01753_));
 INVx1_ASAP7_75t_R _07487_ (.A(_01753_),
    .Y(_01754_));
 INVx1_ASAP7_75t_R _07488_ (.A(_01717_),
    .Y(_01755_));
 NAND2x1_ASAP7_75t_R _07489_ (.A(_01747_),
    .B(_01745_),
    .Y(_01756_));
 AOI21x1_ASAP7_75t_R _07490_ (.A1(net3776),
    .A2(_01755_),
    .B(_01756_),
    .Y(_01757_));
 OAI21x1_ASAP7_75t_R _07491_ (.A1(net3726),
    .A2(_01757_),
    .B(net4172),
    .Y(_01758_));
 AO21x1_ASAP7_75t_R _07492_ (.A1(_01578_),
    .A2(net4385),
    .B(net4342),
    .Y(_01759_));
 NAND2x1_ASAP7_75t_R _07493_ (.A(net4482),
    .B(net4483),
    .Y(_01760_));
 XOR2x2_ASAP7_75t_R _07494_ (.A(_01759_),
    .B(_01760_),
    .Y(_01761_));
 NAND2x1_ASAP7_75t_R _07495_ (.A(net3754),
    .B(net3746),
    .Y(_01762_));
 NOR2x1_ASAP7_75t_R _07496_ (.A(_01761_),
    .B(_01762_),
    .Y(_01763_));
 INVx1_ASAP7_75t_R _07497_ (.A(_01763_),
    .Y(_01764_));
 AOI21x1_ASAP7_75t_R _07498_ (.A1(_01754_),
    .A2(_01758_),
    .B(_01764_),
    .Y(_01765_));
 XOR2x2_ASAP7_75t_R _07499_ (.A(_01683_),
    .B(_01716_),
    .Y(_01766_));
 XOR2x2_ASAP7_75t_R _07500_ (.A(_01717_),
    .B(_01766_),
    .Y(_01767_));
 OAI21x1_ASAP7_75t_R _07501_ (.A1(net3727),
    .A2(_01757_),
    .B(_01767_),
    .Y(_01768_));
 XOR2x2_ASAP7_75t_R _07502_ (.A(net3755),
    .B(_01684_),
    .Y(_01769_));
 NAND3x1_ASAP7_75t_R _07503_ (.A(_01769_),
    .B(_01744_),
    .C(_01739_),
    .Y(_01770_));
 NAND2x2_ASAP7_75t_R _07504_ (.A(_01768_),
    .B(_01770_),
    .Y(_01771_));
 XOR2x2_ASAP7_75t_R _07505_ (.A(_01731_),
    .B(net4049),
    .Y(_01772_));
 NAND3x1_ASAP7_75t_R _07506_ (.A(_01772_),
    .B(_01710_),
    .C(net3775),
    .Y(_01773_));
 OAI21x1_ASAP7_75t_R _07507_ (.A1(_01743_),
    .A2(net3728),
    .B(_01773_),
    .Y(_01774_));
 XOR2x2_ASAP7_75t_R _07508_ (.A(_01774_),
    .B(net3725),
    .Y(_01775_));
 NOR3x1_ASAP7_75t_R _07509_ (.A(_01765_),
    .B(_01771_),
    .C(_01775_),
    .Y(_01776_));
 AOI21x1_ASAP7_75t_R _07510_ (.A1(net3729),
    .A2(net3722),
    .B(net3726),
    .Y(_01777_));
 XOR2x2_ASAP7_75t_R _07511_ (.A(net3741),
    .B(net4098),
    .Y(_01778_));
 AOI21x1_ASAP7_75t_R _07512_ (.A1(_01744_),
    .A2(net5762),
    .B(_01778_),
    .Y(_01779_));
 AOI21x1_ASAP7_75t_R _07513_ (.A1(net3723),
    .A2(_01777_),
    .B(_01779_),
    .Y(_01780_));
 AOI21x1_ASAP7_75t_R _07514_ (.A1(_01744_),
    .A2(net5762),
    .B(net4098),
    .Y(_01781_));
 INVx1_ASAP7_75t_R _07515_ (.A(_01761_),
    .Y(_01782_));
 OAI21x1_ASAP7_75t_R _07516_ (.A1(net3714),
    .A2(_01781_),
    .B(_01782_),
    .Y(_01783_));
 XOR2x2_ASAP7_75t_R _07517_ (.A(_01780_),
    .B(_01783_),
    .Y(_01784_));
 OAI21x1_ASAP7_75t_R _07518_ (.A1(net3676),
    .A2(_01776_),
    .B(_01784_),
    .Y(_01785_));
 NOR2x2_ASAP7_75t_R _07519_ (.A(_01771_),
    .B(_01775_),
    .Y(_01786_));
 NOR3x1_ASAP7_75t_R _07520_ (.A(_01786_),
    .B(_01751_),
    .C(_01780_),
    .Y(_01787_));
 INVx1_ASAP7_75t_R _07521_ (.A(_01787_),
    .Y(_01788_));
 OAI21x1_ASAP7_75t_R _07522_ (.A1(_01781_),
    .A2(_01753_),
    .B(_01763_),
    .Y(_01789_));
 XOR2x2_ASAP7_75t_R _07523_ (.A(net3731),
    .B(_01769_),
    .Y(_01790_));
 NOR2x1_ASAP7_75t_R _07524_ (.A(_01790_),
    .B(_01777_),
    .Y(_01791_));
 AOI211x1_ASAP7_75t_R _07525_ (.A1(net3722),
    .A2(net3729),
    .B(net3742),
    .C(net3727),
    .Y(_01792_));
 NOR2x1_ASAP7_75t_R _07526_ (.A(_01791_),
    .B(_01792_),
    .Y(_01793_));
 AO21x1_ASAP7_75t_R _07527_ (.A1(_01789_),
    .A2(_01751_),
    .B(_01793_),
    .Y(_01794_));
 XNOR2x2_ASAP7_75t_R _07528_ (.A(net3725),
    .B(_01774_),
    .Y(_01795_));
 NOR2x1_ASAP7_75t_R _07529_ (.A(_01771_),
    .B(_01765_),
    .Y(_01796_));
 OAI21x1_ASAP7_75t_R _07530_ (.A1(net3676),
    .A2(net3703),
    .B(_01796_),
    .Y(_01797_));
 NAND2x1_ASAP7_75t_R _07531_ (.A(_01794_),
    .B(_01797_),
    .Y(_01798_));
 AOI21x1_ASAP7_75t_R _07532_ (.A1(_01785_),
    .A2(_01788_),
    .B(_01798_),
    .Y(_01799_));
 NAND2x1_ASAP7_75t_R _07533_ (.A(net3705),
    .B(net3691),
    .Y(_01800_));
 OAI21x1_ASAP7_75t_R _07534_ (.A1(net3677),
    .A2(_01776_),
    .B(net4048),
    .Y(_01801_));
 AOI21x1_ASAP7_75t_R _07535_ (.A1(_01789_),
    .A2(_01786_),
    .B(_01751_),
    .Y(_01802_));
 NAND2x2_ASAP7_75t_R _07536_ (.A(net4023),
    .B(_01802_),
    .Y(_01803_));
 AND2x2_ASAP7_75t_R _07537_ (.A(_01273_),
    .B(net4484),
    .Y(_01804_));
 OAI21x1_ASAP7_75t_R _07538_ (.A1(net4446),
    .A2(net4338),
    .B(net4287),
    .Y(_01805_));
 XNOR2x2_ASAP7_75t_R _07539_ (.A(_01804_),
    .B(_01805_),
    .Y(_01806_));
 AOI21x1_ASAP7_75t_R _07540_ (.A1(_01801_),
    .A2(_01803_),
    .B(net4170),
    .Y(_01807_));
 NAND2x1_ASAP7_75t_R _07541_ (.A(_01807_),
    .B(net3673),
    .Y(_01808_));
 NAND3x1_ASAP7_75t_R _07542_ (.A(_01795_),
    .B(_01793_),
    .C(_01789_),
    .Y(_01809_));
 AO21x1_ASAP7_75t_R _07543_ (.A1(_01796_),
    .A2(_01751_),
    .B(net3703),
    .Y(_01810_));
 NAND2x2_ASAP7_75t_R _07544_ (.A(net5383),
    .B(_01810_),
    .Y(_01811_));
 INVx2_ASAP7_75t_R _07545_ (.A(_01811_),
    .Y(_01812_));
 AOI21x1_ASAP7_75t_R _07546_ (.A1(_01799_),
    .A2(_01808_),
    .B(_01812_),
    .Y(_01813_));
 INVx1_ASAP7_75t_R _07547_ (.A(_01800_),
    .Y(_01814_));
 AOI21x1_ASAP7_75t_R _07548_ (.A1(net3692),
    .A2(_01809_),
    .B(net4023),
    .Y(_01815_));
 AOI211x1_ASAP7_75t_R _07549_ (.A1(net3663),
    .A2(_01789_),
    .B(net3677),
    .C(net4048),
    .Y(_01816_));
 INVx1_ASAP7_75t_R _07550_ (.A(_01806_),
    .Y(_01817_));
 OAI21x1_ASAP7_75t_R _07551_ (.A1(_01816_),
    .A2(_01815_),
    .B(_01817_),
    .Y(_01818_));
 NAND2x1_ASAP7_75t_R _07552_ (.A(_01788_),
    .B(_01785_),
    .Y(_01819_));
 OAI21x1_ASAP7_75t_R _07553_ (.A1(net3662),
    .A2(_01818_),
    .B(_01819_),
    .Y(_01820_));
 AOI211x1_ASAP7_75t_R _07554_ (.A1(net3704),
    .A2(net3692),
    .B(net3675),
    .C(net3674),
    .Y(_01821_));
 INVx1_ASAP7_75t_R _07555_ (.A(_01794_),
    .Y(_01822_));
 NOR2x1_ASAP7_75t_R _07556_ (.A(_01821_),
    .B(_01822_),
    .Y(_01823_));
 XOR2x2_ASAP7_75t_R _07557_ (.A(_01820_),
    .B(net3637),
    .Y(_01824_));
 NAND2x1_ASAP7_75t_R _07558_ (.A(net3637),
    .B(_01813_),
    .Y(_01825_));
 OAI21x1_ASAP7_75t_R _07559_ (.A1(_01813_),
    .A2(_01824_),
    .B(_01825_),
    .Y(_01826_));
 XNOR2x2_ASAP7_75t_R _07560_ (.A(_01783_),
    .B(_01780_),
    .Y(_01827_));
 NOR2x1_ASAP7_75t_R _07561_ (.A(_01827_),
    .B(_01802_),
    .Y(_01828_));
 OAI21x1_ASAP7_75t_R _07562_ (.A1(_01828_),
    .A2(net3652),
    .B(_01823_),
    .Y(_01829_));
 AOI22x1_ASAP7_75t_R _07563_ (.A1(net3618),
    .A2(net3673),
    .B1(_01829_),
    .B2(net3641),
    .Y(_01830_));
 XOR2x2_ASAP7_75t_R _07564_ (.A(_01830_),
    .B(net3616),
    .Y(_01831_));
 OAI21x1_ASAP7_75t_R _07565_ (.A1(net4281),
    .A2(net4229),
    .B(net4290),
    .Y(_01832_));
 XOR2x2_ASAP7_75t_R _07566_ (.A(_01832_),
    .B(net4485),
    .Y(_01833_));
 INVx1_ASAP7_75t_R _07567_ (.A(_01833_),
    .Y(_01834_));
 OAI21x1_ASAP7_75t_R _07568_ (.A1(_01815_),
    .A2(_01816_),
    .B(net3673),
    .Y(_01835_));
 NAND2x1_ASAP7_75t_R _07569_ (.A(_01835_),
    .B(_01799_),
    .Y(_01836_));
 AOI21x1_ASAP7_75t_R _07570_ (.A1(net3641),
    .A2(_01836_),
    .B(net4171),
    .Y(_01837_));
 NAND3x2_ASAP7_75t_R _07571_ (.B(net4171),
    .C(net3641),
    .Y(_01838_),
    .A(net5401));
 INVx2_ASAP7_75t_R _07572_ (.A(_01838_),
    .Y(_01839_));
 NAND2x1_ASAP7_75t_R _07573_ (.A(net3651),
    .B(net3642),
    .Y(_01840_));
 INVx1_ASAP7_75t_R _07574_ (.A(_01840_),
    .Y(_01841_));
 NOR3x1_ASAP7_75t_R _07575_ (.A(_01837_),
    .B(_01839_),
    .C(_01841_),
    .Y(_01842_));
 AO21x1_ASAP7_75t_R _07576_ (.A1(_01809_),
    .A2(net3692),
    .B(_01783_),
    .Y(_01843_));
 OAI21x1_ASAP7_75t_R _07577_ (.A1(net4048),
    .A2(_01802_),
    .B(_01814_),
    .Y(_01844_));
 NAND2x1_ASAP7_75t_R _07578_ (.A(_01843_),
    .B(_01844_),
    .Y(_01845_));
 XOR2x1_ASAP7_75t_R _07579_ (.A(_01845_),
    .Y(_01846_),
    .B(net3618));
 AO211x2_ASAP7_75t_R _07580_ (.A1(net3639),
    .A2(net3619),
    .B(_01845_),
    .C(net3617),
    .Y(_01847_));
 OAI21x1_ASAP7_75t_R _07581_ (.A1(_01813_),
    .A2(_01846_),
    .B(_01847_),
    .Y(_01848_));
 AOI21x1_ASAP7_75t_R _07582_ (.A1(_01842_),
    .A2(net4047),
    .B(_01848_),
    .Y(_01849_));
 OAI21x1_ASAP7_75t_R _07583_ (.A1(net5787),
    .A2(_01826_),
    .B(_01849_),
    .Y(_01850_));
 XNOR2x2_ASAP7_75t_R _07584_ (.A(net3616),
    .B(_01830_),
    .Y(_01851_));
 XOR2x2_ASAP7_75t_R _07585_ (.A(_01850_),
    .B(net3595),
    .Y(_01852_));
 NAND2x1_ASAP7_75t_R _07586_ (.A(net4338),
    .B(net4290),
    .Y(_01853_));
 NOR2x1_ASAP7_75t_R _07587_ (.A(net4487),
    .B(net4486),
    .Y(_01854_));
 INVx1_ASAP7_75t_R _07588_ (.A(_01854_),
    .Y(_01855_));
 XOR2x2_ASAP7_75t_R _07589_ (.A(_01853_),
    .B(_01855_),
    .Y(_01856_));
 INVx1_ASAP7_75t_R _07590_ (.A(_01856_),
    .Y(_01857_));
 OAI21x1_ASAP7_75t_R _07591_ (.A1(net3662),
    .A2(net3638),
    .B(net3619),
    .Y(_01858_));
 NAND2x1_ASAP7_75t_R _07592_ (.A(net3640),
    .B(_01858_),
    .Y(_01859_));
 INVx1_ASAP7_75t_R _07593_ (.A(_01846_),
    .Y(_01860_));
 AOI211x1_ASAP7_75t_R _07594_ (.A1(net3619),
    .A2(net3638),
    .B(net3617),
    .C(net3614),
    .Y(_01861_));
 AOI21x1_ASAP7_75t_R _07595_ (.A1(_01859_),
    .A2(_01860_),
    .B(_01861_),
    .Y(_01862_));
 NAND2x1p5_ASAP7_75t_R _07596_ (.A(_01831_),
    .B(_01862_),
    .Y(_01863_));
 AOI21x1_ASAP7_75t_R _07597_ (.A1(net3651),
    .A2(net3642),
    .B(net3662),
    .Y(_01864_));
 NOR2x1_ASAP7_75t_R _07598_ (.A(_01829_),
    .B(_01864_),
    .Y(_01865_));
 OAI21x1_ASAP7_75t_R _07599_ (.A1(_01812_),
    .A2(_01865_),
    .B(net4097),
    .Y(_01866_));
 NAND3x1_ASAP7_75t_R _07600_ (.A(_01866_),
    .B(_01840_),
    .C(_01838_),
    .Y(_01867_));
 NOR2x1_ASAP7_75t_R _07601_ (.A(net4096),
    .B(_01867_),
    .Y(_01868_));
 INVx2_ASAP7_75t_R _07602_ (.A(_01826_),
    .Y(_01869_));
 OAI21x1_ASAP7_75t_R _07603_ (.A1(net3565),
    .A2(_01868_),
    .B(_01869_),
    .Y(_01870_));
 NOR2x1_ASAP7_75t_R _07604_ (.A(net4047),
    .B(_01870_),
    .Y(_01871_));
 NOR2x2_ASAP7_75t_R _07605_ (.A(_01839_),
    .B(net3596),
    .Y(_01872_));
 INVx1_ASAP7_75t_R _07606_ (.A(net3580),
    .Y(_01873_));
 NAND3x1_ASAP7_75t_R _07607_ (.A(net3581),
    .B(net3582),
    .C(net3597),
    .Y(_01874_));
 AOI21x1_ASAP7_75t_R _07608_ (.A1(net3553),
    .A2(_01874_),
    .B(net4096),
    .Y(_01875_));
 NOR3x1_ASAP7_75t_R _07609_ (.A(_01871_),
    .B(_01873_),
    .C(_01875_),
    .Y(_01876_));
 AND3x1_ASAP7_75t_R _07610_ (.A(_01866_),
    .B(_01834_),
    .C(_01838_),
    .Y(_01877_));
 AND3x1_ASAP7_75t_R _07611_ (.A(_01877_),
    .B(_01826_),
    .C(net3615),
    .Y(_01878_));
 XOR2x2_ASAP7_75t_R _07612_ (.A(net3596),
    .B(net3615),
    .Y(_01879_));
 AOI21x1_ASAP7_75t_R _07613_ (.A1(net3579),
    .A2(_01870_),
    .B(net3578),
    .Y(_01880_));
 OAI21x1_ASAP7_75t_R _07614_ (.A1(_01869_),
    .A2(_01868_),
    .B(net3583),
    .Y(_01881_));
 NAND2x2_ASAP7_75t_R _07615_ (.A(_01881_),
    .B(_01850_),
    .Y(_01882_));
 INVx1_ASAP7_75t_R _07616_ (.A(_01882_),
    .Y(_01883_));
 OAI21x1_ASAP7_75t_R _07617_ (.A1(net3552),
    .A2(_01880_),
    .B(_01883_),
    .Y(_01884_));
 AOI21x1_ASAP7_75t_R _07618_ (.A1(_01857_),
    .A2(_01876_),
    .B(_01884_),
    .Y(_01885_));
 OAI21x1_ASAP7_75t_R _07619_ (.A1(net3541),
    .A2(_01885_),
    .B(net4095),
    .Y(_01886_));
 NOR2x1_ASAP7_75t_R _07620_ (.A(_01851_),
    .B(_01848_),
    .Y(_01887_));
 NAND3x1_ASAP7_75t_R _07621_ (.A(_01872_),
    .B(net4047),
    .C(net3615),
    .Y(_01888_));
 AOI21x1_ASAP7_75t_R _07622_ (.A1(_01887_),
    .A2(_01888_),
    .B(_01826_),
    .Y(_01889_));
 NAND2x2_ASAP7_75t_R _07623_ (.A(_01889_),
    .B(net4096),
    .Y(_01890_));
 NOR2x1_ASAP7_75t_R _07624_ (.A(net3584),
    .B(_01863_),
    .Y(_01891_));
 OAI21x1_ASAP7_75t_R _07625_ (.A1(_01891_),
    .A2(net3566),
    .B(net4047),
    .Y(_01892_));
 NAND3x2_ASAP7_75t_R _07626_ (.B(_01892_),
    .C(_01890_),
    .Y(_01893_),
    .A(net3580));
 INVx1_ASAP7_75t_R _07627_ (.A(_01878_),
    .Y(_01894_));
 INVx1_ASAP7_75t_R _07628_ (.A(net3579),
    .Y(_01895_));
 INVx1_ASAP7_75t_R _07629_ (.A(_01879_),
    .Y(_01896_));
 OAI21x1_ASAP7_75t_R _07630_ (.A1(_01895_),
    .A2(_01889_),
    .B(_01896_),
    .Y(_01897_));
 AOI21x1_ASAP7_75t_R _07631_ (.A1(_01894_),
    .A2(_01897_),
    .B(_01882_),
    .Y(_01898_));
 OAI21x1_ASAP7_75t_R _07632_ (.A1(net4168),
    .A2(_01893_),
    .B(_01898_),
    .Y(_01899_));
 INVx3_ASAP7_75t_R _07633_ (.A(_01852_),
    .Y(_01900_));
 NAND3x2_ASAP7_75t_R _07634_ (.B(net4169),
    .C(_01900_),
    .Y(_01901_),
    .A(net5389));
 NAND2x2_ASAP7_75t_R _07635_ (.A(_01886_),
    .B(_01901_),
    .Y(_01902_));
 INVx1_ASAP7_75t_R _07636_ (.A(net3464),
    .Y(_01903_));
 NAND2x2_ASAP7_75t_R _07637_ (.A(_01900_),
    .B(net5390),
    .Y(_01904_));
 NAND2x2_ASAP7_75t_R _07638_ (.A(net3538),
    .B(net3537),
    .Y(_01905_));
 OAI21x1_ASAP7_75t_R _07639_ (.A1(net4169),
    .A2(net3521),
    .B(_01905_),
    .Y(_01906_));
 XOR2x2_ASAP7_75t_R _07640_ (.A(_01906_),
    .B(net3522),
    .Y(_01907_));
 NOR2x1p5_ASAP7_75t_R _07641_ (.A(net3522),
    .B(_01904_),
    .Y(_01908_));
 AOI21x1_ASAP7_75t_R _07642_ (.A1(_01904_),
    .A2(_01907_),
    .B(_01908_),
    .Y(_01909_));
 AO21x1_ASAP7_75t_R _07643_ (.A1(_01576_),
    .A2(net4387),
    .B(net4342),
    .Y(_01910_));
 XOR2x2_ASAP7_75t_R _07644_ (.A(_01910_),
    .B(net4386),
    .Y(_01911_));
 NAND2x1_ASAP7_75t_R _07645_ (.A(net5822),
    .B(net3540),
    .Y(_01912_));
 INVx1_ASAP7_75t_R _07646_ (.A(_01912_),
    .Y(_01913_));
 NAND3x1_ASAP7_75t_R _07647_ (.A(_01901_),
    .B(_01886_),
    .C(_01913_),
    .Y(_01914_));
 NAND3x1_ASAP7_75t_R _07648_ (.A(net3540),
    .B(net3539),
    .C(_01857_),
    .Y(_01915_));
 XOR2x2_ASAP7_75t_R _07649_ (.A(_01875_),
    .B(net3580),
    .Y(_01916_));
 XOR2x2_ASAP7_75t_R _07650_ (.A(_01915_),
    .B(_01916_),
    .Y(_01917_));
 OAI21x1_ASAP7_75t_R _07651_ (.A1(net5456),
    .A2(net3485),
    .B(_01917_),
    .Y(_01918_));
 INVx1_ASAP7_75t_R _07652_ (.A(_01916_),
    .Y(_01919_));
 NAND3x1_ASAP7_75t_R _07653_ (.A(net5389),
    .B(_01919_),
    .C(_01900_),
    .Y(_01920_));
 INVx1_ASAP7_75t_R _07654_ (.A(_01905_),
    .Y(_01921_));
 AOI22x1_ASAP7_75t_R _07655_ (.A1(net3492),
    .A2(_01900_),
    .B1(net3506),
    .B2(net4095),
    .Y(_01922_));
 NAND2x1_ASAP7_75t_R _07656_ (.A(_01921_),
    .B(_01922_),
    .Y(_01923_));
 OAI22x1_ASAP7_75t_R _07657_ (.A1(net3521),
    .A2(net4169),
    .B1(net3505),
    .B2(net3541),
    .Y(_01924_));
 NAND2x1_ASAP7_75t_R _07658_ (.A(net3519),
    .B(_01924_),
    .Y(_01925_));
 AOI22x1_ASAP7_75t_R _07659_ (.A1(_01920_),
    .A2(_01918_),
    .B1(_01923_),
    .B2(_01925_),
    .Y(_01926_));
 OAI21x1_ASAP7_75t_R _07660_ (.A1(net4166),
    .A2(_01914_),
    .B(_01926_),
    .Y(_01927_));
 NAND2x1_ASAP7_75t_R _07661_ (.A(net3463),
    .B(net3449),
    .Y(_01928_));
 XOR2x2_ASAP7_75t_R _07662_ (.A(net3464),
    .B(net4167),
    .Y(_01929_));
 AO21x1_ASAP7_75t_R _07663_ (.A1(net3449),
    .A2(net3463),
    .B(_01929_),
    .Y(_01930_));
 OAI21x1_ASAP7_75t_R _07664_ (.A1(_01903_),
    .A2(_01928_),
    .B(_01930_),
    .Y(_01931_));
 INVx3_ASAP7_75t_R _07665_ (.A(_01909_),
    .Y(_01932_));
 AOI211x1_ASAP7_75t_R _07666_ (.A1(_01926_),
    .A2(_01914_),
    .B(net4167),
    .C(_01932_),
    .Y(_01933_));
 INVx1_ASAP7_75t_R _07667_ (.A(_01911_),
    .Y(_01934_));
 AOI21x1_ASAP7_75t_R _07668_ (.A1(_01927_),
    .A2(net5388),
    .B(net4094),
    .Y(_01935_));
 NAND2x1_ASAP7_75t_R _07669_ (.A(net4287),
    .B(net4382),
    .Y(_01936_));
 XNOR2x2_ASAP7_75t_R _07670_ (.A(net4439),
    .B(_01936_),
    .Y(_01937_));
 INVx1_ASAP7_75t_R _07671_ (.A(_01937_),
    .Y(_01938_));
 OAI21x1_ASAP7_75t_R _07672_ (.A1(_01935_),
    .A2(_01933_),
    .B(_01938_),
    .Y(_01939_));
 XOR2x2_ASAP7_75t_R _07673_ (.A(_01931_),
    .B(net3417),
    .Y(_01940_));
 NOR2x2_ASAP7_75t_R _07674_ (.A(_01939_),
    .B(net3464),
    .Y(_01941_));
 AOI21x1_ASAP7_75t_R _07675_ (.A1(net3520),
    .A2(net3491),
    .B(net4169),
    .Y(_01942_));
 XOR2x2_ASAP7_75t_R _07676_ (.A(_01942_),
    .B(net3518),
    .Y(_01943_));
 INVx1_ASAP7_75t_R _07677_ (.A(_01943_),
    .Y(_01944_));
 NAND3x1_ASAP7_75t_R _07678_ (.A(net3484),
    .B(net3476),
    .C(_01934_),
    .Y(_01945_));
 AOI21x1_ASAP7_75t_R _07679_ (.A1(_01909_),
    .A2(_01927_),
    .B(_01945_),
    .Y(_01946_));
 OR3x1_ASAP7_75t_R _07680_ (.A(_01945_),
    .B(_01909_),
    .C(net3518),
    .Y(_01947_));
 OAI21x1_ASAP7_75t_R _07681_ (.A1(_01944_),
    .A2(_01946_),
    .B(_01947_),
    .Y(_01948_));
 INVx1_ASAP7_75t_R _07682_ (.A(_01920_),
    .Y(_01949_));
 INVx2_ASAP7_75t_R _07683_ (.A(_01918_),
    .Y(_01950_));
 NOR2x1_ASAP7_75t_R _07684_ (.A(_01949_),
    .B(_01950_),
    .Y(_01951_));
 XOR2x2_ASAP7_75t_R _07685_ (.A(_01921_),
    .B(_01924_),
    .Y(_01952_));
 OAI21x1_ASAP7_75t_R _07686_ (.A1(_01950_),
    .A2(_01949_),
    .B(_01952_),
    .Y(_01953_));
 NOR2x1_ASAP7_75t_R _07687_ (.A(net3518),
    .B(_01902_),
    .Y(_01954_));
 AOI22x1_ASAP7_75t_R _07688_ (.A1(_01909_),
    .A2(_01953_),
    .B1(_01954_),
    .B2(net4094),
    .Y(_01955_));
 XNOR2x2_ASAP7_75t_R _07689_ (.A(_01951_),
    .B(_01955_),
    .Y(_01956_));
 NAND2x2_ASAP7_75t_R _07690_ (.A(_01956_),
    .B(_01948_),
    .Y(_01957_));
 INVx1_ASAP7_75t_R _07691_ (.A(_01952_),
    .Y(_01958_));
 AOI21x1_ASAP7_75t_R _07692_ (.A1(net4094),
    .A2(net3444),
    .B(_01951_),
    .Y(_01959_));
 NAND3x1_ASAP7_75t_R _07693_ (.A(_01959_),
    .B(net5424),
    .C(_01958_),
    .Y(_01960_));
 OAI21x1_ASAP7_75t_R _07694_ (.A1(net3475),
    .A2(net3427),
    .B(_01960_),
    .Y(_01961_));
 INVx2_ASAP7_75t_R _07695_ (.A(_01961_),
    .Y(_01962_));
 OAI21x1_ASAP7_75t_R _07696_ (.A1(_01957_),
    .A2(_01941_),
    .B(_01962_),
    .Y(_01963_));
 NAND2x1_ASAP7_75t_R _07697_ (.A(_01940_),
    .B(net3377),
    .Y(_01964_));
 INVx1_ASAP7_75t_R _07698_ (.A(_01931_),
    .Y(_01965_));
 XOR2x2_ASAP7_75t_R _07699_ (.A(net5450),
    .B(net3446),
    .Y(_01966_));
 AOI21x1_ASAP7_75t_R _07700_ (.A1(net4094),
    .A2(net3444),
    .B(net3445),
    .Y(_01967_));
 XOR2x2_ASAP7_75t_R _07701_ (.A(_01945_),
    .B(_01943_),
    .Y(_01968_));
 OAI21x1_ASAP7_75t_R _07702_ (.A1(net3447),
    .A2(_01967_),
    .B(_01968_),
    .Y(_01969_));
 NAND3x1_ASAP7_75t_R _07703_ (.A(net3449),
    .B(net3463),
    .C(_01944_),
    .Y(_01970_));
 NAND2x1_ASAP7_75t_R _07704_ (.A(_01969_),
    .B(_01970_),
    .Y(_01971_));
 NOR2x1_ASAP7_75t_R _07705_ (.A(_01966_),
    .B(_01971_),
    .Y(_01972_));
 OAI21x1_ASAP7_75t_R _07706_ (.A1(net3448),
    .A2(_01967_),
    .B(net4167),
    .Y(_01973_));
 INVx1_ASAP7_75t_R _07707_ (.A(net3430),
    .Y(_01974_));
 AOI21x1_ASAP7_75t_R _07708_ (.A1(_01973_),
    .A2(_01974_),
    .B(net4165),
    .Y(_01975_));
 NAND2x1_ASAP7_75t_R _07709_ (.A(net3450),
    .B(_01975_),
    .Y(_01976_));
 AOI21x1_ASAP7_75t_R _07710_ (.A1(_01972_),
    .A2(_01976_),
    .B(net3403),
    .Y(_01977_));
 NAND2x1_ASAP7_75t_R _07711_ (.A(_01965_),
    .B(_01977_),
    .Y(_01978_));
 NAND2x1_ASAP7_75t_R _07712_ (.A(_01978_),
    .B(_01964_),
    .Y(_01979_));
 NOR2x2_ASAP7_75t_R _07713_ (.A(_01963_),
    .B(net4093),
    .Y(_01980_));
 OAI21x1_ASAP7_75t_R _07714_ (.A1(net3430),
    .A2(net3429),
    .B(_01903_),
    .Y(_01981_));
 NAND3x1_ASAP7_75t_R _07715_ (.A(net3415),
    .B(net3416),
    .C(_01981_),
    .Y(_01982_));
 AOI21x1_ASAP7_75t_R _07716_ (.A1(_01982_),
    .A2(net3392),
    .B(net4165),
    .Y(_01983_));
 NOR2x1_ASAP7_75t_R _07717_ (.A(net4342),
    .B(_01576_),
    .Y(_01984_));
 XOR2x2_ASAP7_75t_R _07718_ (.A(_01984_),
    .B(net4440),
    .Y(_01985_));
 NAND2x1_ASAP7_75t_R _07719_ (.A(_01973_),
    .B(_01974_),
    .Y(_01986_));
 INVx1_ASAP7_75t_R _07720_ (.A(_01986_),
    .Y(_01987_));
 NOR2x1_ASAP7_75t_R _07721_ (.A(_01985_),
    .B(_01987_),
    .Y(_01988_));
 INVx1_ASAP7_75t_R _07722_ (.A(_01988_),
    .Y(_01989_));
 NOR3x2_ASAP7_75t_R _07723_ (.B(_01980_),
    .C(_01989_),
    .Y(_01990_),
    .A(_01983_));
 NOR2x1_ASAP7_75t_R _07724_ (.A(net3355),
    .B(_01990_),
    .Y(_01991_));
 INVx1_ASAP7_75t_R _07725_ (.A(_01991_),
    .Y(_01992_));
 NOR2x2_ASAP7_75t_R _07726_ (.A(_01980_),
    .B(_01983_),
    .Y(_01993_));
 NAND2x1_ASAP7_75t_R _07727_ (.A(net3375),
    .B(_01993_),
    .Y(_01994_));
 XOR2x2_ASAP7_75t_R _07728_ (.A(net3405),
    .B(net3402),
    .Y(_01995_));
 NOR2x1_ASAP7_75t_R _07729_ (.A(net5819),
    .B(net3403),
    .Y(_01996_));
 INVx1_ASAP7_75t_R _07730_ (.A(_01996_),
    .Y(_01997_));
 OAI21x1_ASAP7_75t_R _07731_ (.A1(net3376),
    .A2(_01995_),
    .B(_01997_),
    .Y(_01998_));
 NOR2x1_ASAP7_75t_R _07732_ (.A(_01998_),
    .B(_01979_),
    .Y(_01999_));
 OAI21x1_ASAP7_75t_R _07733_ (.A1(net3464),
    .A2(net3418),
    .B(net5820),
    .Y(_02000_));
 AO21x1_ASAP7_75t_R _07734_ (.A1(_02000_),
    .A2(net3414),
    .B(net3392),
    .Y(_02001_));
 OA21x2_ASAP7_75t_R _07735_ (.A1(net3414),
    .A2(net3378),
    .B(_02001_),
    .Y(_02002_));
 INVx2_ASAP7_75t_R _07736_ (.A(_02002_),
    .Y(_02003_));
 AOI21x1_ASAP7_75t_R _07737_ (.A1(_01994_),
    .A2(_01999_),
    .B(_02003_),
    .Y(_02004_));
 OA21x2_ASAP7_75t_R _07738_ (.A1(net3354),
    .A2(net3367),
    .B(net3355),
    .Y(_02005_));
 INVx1_ASAP7_75t_R _07739_ (.A(_02005_),
    .Y(_02006_));
 OAI21x1_ASAP7_75t_R _07740_ (.A1(_01992_),
    .A2(_02004_),
    .B(_02006_),
    .Y(_02007_));
 XOR2x2_ASAP7_75t_R _07741_ (.A(net5770),
    .B(net3416),
    .Y(_02008_));
 AOI21x1_ASAP7_75t_R _07742_ (.A1(net3377),
    .A2(_02008_),
    .B(_01996_),
    .Y(_02009_));
 OA21x2_ASAP7_75t_R _07743_ (.A1(net3392),
    .A2(net3418),
    .B(_01965_),
    .Y(_02010_));
 AOI211x1_ASAP7_75t_R _07744_ (.A1(net3404),
    .A2(net3392),
    .B(net3418),
    .C(_01965_),
    .Y(_02011_));
 NOR2x1_ASAP7_75t_R _07745_ (.A(_02010_),
    .B(_02011_),
    .Y(_02012_));
 NAND2x1_ASAP7_75t_R _07746_ (.A(_02012_),
    .B(_02009_),
    .Y(_02013_));
 OAI21x1_ASAP7_75t_R _07747_ (.A1(_02013_),
    .A2(_01990_),
    .B(_02002_),
    .Y(_02014_));
 NOR3x1_ASAP7_75t_R _07748_ (.A(_01980_),
    .B(_01983_),
    .C(net4164),
    .Y(_02015_));
 XOR2x2_ASAP7_75t_R _07749_ (.A(net3401),
    .B(net4093),
    .Y(_02016_));
 NOR2x1_ASAP7_75t_R _07750_ (.A(net3391),
    .B(net3378),
    .Y(_02017_));
 AOI21x1_ASAP7_75t_R _07751_ (.A1(net3378),
    .A2(_02016_),
    .B(_02017_),
    .Y(_02018_));
 XOR2x2_ASAP7_75t_R _07752_ (.A(_02015_),
    .B(_02018_),
    .Y(_02019_));
 INVx1_ASAP7_75t_R _07753_ (.A(_02018_),
    .Y(_02020_));
 NOR3x1_ASAP7_75t_R _07754_ (.A(net5444),
    .B(_02020_),
    .C(_02003_),
    .Y(_02021_));
 AOI21x1_ASAP7_75t_R _07755_ (.A1(net5439),
    .A2(_02019_),
    .B(_02021_),
    .Y(_02022_));
 NOR2x1p5_ASAP7_75t_R _07756_ (.A(_02007_),
    .B(_02022_),
    .Y(_02023_));
 NOR2x1_ASAP7_75t_R _07757_ (.A(net3354),
    .B(net3352),
    .Y(_02024_));
 INVx1_ASAP7_75t_R _07758_ (.A(_02024_),
    .Y(_02025_));
 AO21x1_ASAP7_75t_R _07759_ (.A1(_01991_),
    .A2(_02003_),
    .B(net3366),
    .Y(_02026_));
 NAND2x1p5_ASAP7_75t_R _07760_ (.A(_02025_),
    .B(_02026_),
    .Y(_02027_));
 INVx2_ASAP7_75t_R _07761_ (.A(_02027_),
    .Y(_02028_));
 INVx1_ASAP7_75t_R _07762_ (.A(net4164),
    .Y(_02029_));
 XOR2x2_ASAP7_75t_R _07763_ (.A(_02029_),
    .B(net5439),
    .Y(_02030_));
 NAND2x2_ASAP7_75t_R _07764_ (.A(net3353),
    .B(_02030_),
    .Y(_02031_));
 AND5x1_ASAP7_75t_R _07765_ (.A(net4595),
    .B(net4390),
    .C(_01152_),
    .D(net4537),
    .E(net4538),
    .Y(_02032_));
 BUFx3_ASAP7_75t_R place3022 (.A(_05129_),
    .Y(net3022));
 AO21x1_ASAP7_75t_R _07767_ (.A1(_02032_),
    .A2(net4531),
    .B(net4342),
    .Y(_02034_));
 NAND2x1_ASAP7_75t_R _07768_ (.A(net4437),
    .B(net4476),
    .Y(_02035_));
 XOR2x2_ASAP7_75t_R _07769_ (.A(_02034_),
    .B(_02035_),
    .Y(_02036_));
 OAI22x1_ASAP7_75t_R _07770_ (.A1(_02023_),
    .A2(_02028_),
    .B1(_02031_),
    .B2(net4227),
    .Y(_02037_));
 XOR2x2_ASAP7_75t_R _07771_ (.A(net3267),
    .B(net3300),
    .Y(_02038_));
 XOR2x2_ASAP7_75t_R _07772_ (.A(net4164),
    .B(net5439),
    .Y(_02039_));
 NOR2x2_ASAP7_75t_R _07773_ (.A(_02036_),
    .B(_02039_),
    .Y(_02040_));
 INVx1_ASAP7_75t_R _07774_ (.A(_02040_),
    .Y(_02041_));
 AOI21x1_ASAP7_75t_R _07775_ (.A1(net3338),
    .A2(net5439),
    .B(net3337),
    .Y(_02042_));
 NOR2x1_ASAP7_75t_R _07776_ (.A(net3353),
    .B(net5439),
    .Y(_02043_));
 XOR2x2_ASAP7_75t_R _07777_ (.A(_01993_),
    .B(net4164),
    .Y(_02044_));
 INVx1_ASAP7_75t_R _07778_ (.A(_02044_),
    .Y(_02045_));
 NOR2x1_ASAP7_75t_R _07779_ (.A(_02004_),
    .B(_02045_),
    .Y(_02046_));
 NOR2x1_ASAP7_75t_R _07780_ (.A(_02046_),
    .B(_02043_),
    .Y(_02047_));
 NOR2x1_ASAP7_75t_R _07781_ (.A(net3300),
    .B(_02047_),
    .Y(_02048_));
 AOI21x1_ASAP7_75t_R _07782_ (.A1(net3317),
    .A2(_02048_),
    .B(net3280),
    .Y(_02049_));
 OAI21x1_ASAP7_75t_R _07783_ (.A1(_02041_),
    .A2(_02049_),
    .B(net3279),
    .Y(_02050_));
 XOR2x2_ASAP7_75t_R _07784_ (.A(net3351),
    .B(_02020_),
    .Y(_02051_));
 NAND3x1_ASAP7_75t_R _07785_ (.A(net3352),
    .B(net3350),
    .C(net3367),
    .Y(_02052_));
 OAI21x1_ASAP7_75t_R _07786_ (.A1(net3321),
    .A2(_02051_),
    .B(_02052_),
    .Y(_02053_));
 OAI21x1_ASAP7_75t_R _07787_ (.A1(net3297),
    .A2(net3316),
    .B(_02053_),
    .Y(_02054_));
 OAI21x1_ASAP7_75t_R _07788_ (.A1(net3301),
    .A2(_02054_),
    .B(net3299),
    .Y(_02055_));
 NAND2x1_ASAP7_75t_R _07789_ (.A(net3336),
    .B(net5439),
    .Y(_02056_));
 INVx1_ASAP7_75t_R _07790_ (.A(net3353),
    .Y(_02057_));
 NAND2x1_ASAP7_75t_R _07791_ (.A(_02057_),
    .B(net3322),
    .Y(_02058_));
 NAND2x2_ASAP7_75t_R _07792_ (.A(_02058_),
    .B(_02056_),
    .Y(_02059_));
 NAND3x1_ASAP7_75t_R _07793_ (.A(_02055_),
    .B(_02040_),
    .C(_02059_),
    .Y(_02060_));
 NAND2x1_ASAP7_75t_R _07794_ (.A(_02050_),
    .B(_02060_),
    .Y(_02061_));
 NAND2x1_ASAP7_75t_R _07795_ (.A(net4287),
    .B(net4331),
    .Y(_02062_));
 INVx1_ASAP7_75t_R _07796_ (.A(net4436),
    .Y(_02063_));
 XOR2x2_ASAP7_75t_R _07797_ (.A(_02062_),
    .B(_02063_),
    .Y(_02064_));
 AOI21x1_ASAP7_75t_R _07798_ (.A1(_02023_),
    .A2(_02031_),
    .B(_02028_),
    .Y(_02065_));
 NOR2x1_ASAP7_75t_R _07799_ (.A(_02057_),
    .B(_02039_),
    .Y(_02066_));
 NAND2x1_ASAP7_75t_R _07800_ (.A(_02066_),
    .B(_02023_),
    .Y(_02067_));
 NAND3x1_ASAP7_75t_R _07801_ (.A(_02065_),
    .B(net4227),
    .C(_02067_),
    .Y(_02068_));
 NOR2x2_ASAP7_75t_R _07802_ (.A(_02065_),
    .B(net4228),
    .Y(_02069_));
 INVx3_ASAP7_75t_R _07803_ (.A(_02069_),
    .Y(_02070_));
 NAND3x2_ASAP7_75t_R _07804_ (.B(net3320),
    .C(_02068_),
    .Y(_02071_),
    .A(_02070_));
 NOR2x2_ASAP7_75t_R _07805_ (.A(net4162),
    .B(_02071_),
    .Y(_02072_));
 NOR2x1p5_ASAP7_75t_R _07806_ (.A(net3223),
    .B(_02072_),
    .Y(_02073_));
 AOI221x1_ASAP7_75t_R _07807_ (.A1(net3301),
    .A2(net3299),
    .B1(_02047_),
    .B2(_02040_),
    .C(net3300),
    .Y(_02074_));
 XOR2x2_ASAP7_75t_R _07808_ (.A(_02074_),
    .B(net3318),
    .Y(_02075_));
 AOI21x1_ASAP7_75t_R _07809_ (.A1(net3245),
    .A2(_02073_),
    .B(net3250),
    .Y(_02076_));
 AOI21x1_ASAP7_75t_R _07810_ (.A1(net3250),
    .A2(_02073_),
    .B(_02076_),
    .Y(_02077_));
 INVx2_ASAP7_75t_R _07811_ (.A(_02077_),
    .Y(_02078_));
 NAND3x1_ASAP7_75t_R _07812_ (.A(_02059_),
    .B(net3317),
    .C(net5765),
    .Y(_02079_));
 AOI21x1_ASAP7_75t_R _07813_ (.A1(net3299),
    .A2(_02079_),
    .B(_02041_),
    .Y(_02080_));
 XOR2x2_ASAP7_75t_R _07814_ (.A(_02080_),
    .B(net3278),
    .Y(_02081_));
 XOR2x2_ASAP7_75t_R _07815_ (.A(_02037_),
    .B(net3296),
    .Y(_02082_));
 NOR2x1p5_ASAP7_75t_R _07816_ (.A(_02061_),
    .B(_02082_),
    .Y(_02083_));
 OAI22x1_ASAP7_75t_R _07817_ (.A1(net5441),
    .A2(net3245),
    .B1(net4162),
    .B2(net3222),
    .Y(_02084_));
 NOR2x1_ASAP7_75t_R _07818_ (.A(net3236),
    .B(_02084_),
    .Y(_02085_));
 NAND2x1_ASAP7_75t_R _07819_ (.A(net3236),
    .B(_02084_),
    .Y(_02086_));
 INVx1_ASAP7_75t_R _07820_ (.A(_02086_),
    .Y(_02087_));
 INVx1_ASAP7_75t_R _07821_ (.A(net4228),
    .Y(_02088_));
 NAND2x1_ASAP7_75t_R _07822_ (.A(net5765),
    .B(_02042_),
    .Y(_02089_));
 OAI21x1_ASAP7_75t_R _07823_ (.A1(_02089_),
    .A2(net3295),
    .B(net3299),
    .Y(_02090_));
 AOI21x1_ASAP7_75t_R _07824_ (.A1(_02088_),
    .A2(_02090_),
    .B(net3320),
    .Y(_02091_));
 NOR2x1_ASAP7_75t_R _07825_ (.A(_02080_),
    .B(_02091_),
    .Y(_02092_));
 INVx1_ASAP7_75t_R _07826_ (.A(_02075_),
    .Y(_02093_));
 INVx1_ASAP7_75t_R _07827_ (.A(_02092_),
    .Y(_02094_));
 NAND3x1_ASAP7_75t_R _07828_ (.A(_02081_),
    .B(_02094_),
    .C(_02038_),
    .Y(_02095_));
 NAND2x2_ASAP7_75t_R _07829_ (.A(net5454),
    .B(net3249),
    .Y(_02096_));
 NOR2x1_ASAP7_75t_R _07830_ (.A(_02064_),
    .B(_02096_),
    .Y(_02097_));
 INVx1_ASAP7_75t_R _07831_ (.A(_02097_),
    .Y(_02098_));
 AOI21x1_ASAP7_75t_R _07832_ (.A1(_02093_),
    .A2(_02095_),
    .B(_02098_),
    .Y(_02099_));
 NAND2x1_ASAP7_75t_R _07833_ (.A(net3246),
    .B(_02072_),
    .Y(_02100_));
 OAI21x1_ASAP7_75t_R _07834_ (.A1(net3235),
    .A2(_02099_),
    .B(_02100_),
    .Y(_02101_));
 OAI21x1_ASAP7_75t_R _07835_ (.A1(_02085_),
    .A2(_02087_),
    .B(_02101_),
    .Y(_02102_));
 NAND2x1_ASAP7_75t_R _07836_ (.A(net4378),
    .B(net4287),
    .Y(_02103_));
 INVx1_ASAP7_75t_R _07837_ (.A(net4480),
    .Y(_02104_));
 INVx1_ASAP7_75t_R _07838_ (.A(net4532),
    .Y(_02105_));
 NAND2x1_ASAP7_75t_R _07839_ (.A(_02104_),
    .B(_02105_),
    .Y(_02106_));
 XOR2x2_ASAP7_75t_R _07840_ (.A(_02103_),
    .B(_02106_),
    .Y(_02107_));
 AOI211x1_ASAP7_75t_R _07841_ (.A1(_02071_),
    .A2(_02083_),
    .B(net3246),
    .C(net4162),
    .Y(_02108_));
 OAI21x1_ASAP7_75t_R _07842_ (.A1(net4162),
    .A2(net5392),
    .B(net5440),
    .Y(_02109_));
 INVx1_ASAP7_75t_R _07843_ (.A(net4162),
    .Y(_02110_));
 AOI21x1_ASAP7_75t_R _07844_ (.A1(_02093_),
    .A2(_02109_),
    .B(_02110_),
    .Y(_02111_));
 INVx1_ASAP7_75t_R _07845_ (.A(net3220),
    .Y(_02112_));
 OAI21x1_ASAP7_75t_R _07846_ (.A1(_02111_),
    .A2(_02108_),
    .B(_02112_),
    .Y(_02113_));
 NOR2x1_ASAP7_75t_R _07847_ (.A(net4159),
    .B(_02113_),
    .Y(_02114_));
 NOR3x1_ASAP7_75t_R _07848_ (.A(net3223),
    .B(net3244),
    .C(net3235),
    .Y(_02115_));
 OAI21x1_ASAP7_75t_R _07849_ (.A1(net3247),
    .A2(_02115_),
    .B(net3206),
    .Y(_02116_));
 NOR2x1_ASAP7_75t_R _07850_ (.A(net3277),
    .B(net3298),
    .Y(_02117_));
 NOR3x1_ASAP7_75t_R _07851_ (.A(net3266),
    .B(_02117_),
    .C(net4161),
    .Y(_02118_));
 NOR3x1_ASAP7_75t_R _07852_ (.A(_02118_),
    .B(net3319),
    .C(net3248),
    .Y(_02119_));
 AND3x1_ASAP7_75t_R _07853_ (.A(_02119_),
    .B(_02110_),
    .C(net3246),
    .Y(_02120_));
 AOI21x1_ASAP7_75t_R _07854_ (.A1(net3221),
    .A2(_02116_),
    .B(_02120_),
    .Y(_02121_));
 AOI211x1_ASAP7_75t_R _07855_ (.A1(_02078_),
    .A2(_02102_),
    .B(net3157),
    .C(net3182),
    .Y(_02122_));
 INVx1_ASAP7_75t_R _07856_ (.A(_02085_),
    .Y(_02123_));
 NAND2x1_ASAP7_75t_R _07857_ (.A(net3184),
    .B(net3171),
    .Y(_02124_));
 XOR2x2_ASAP7_75t_R _07858_ (.A(_02122_),
    .B(_02124_),
    .Y(_02125_));
 NAND2x2_ASAP7_75t_R _07859_ (.A(_02038_),
    .B(_02081_),
    .Y(_02126_));
 NOR2x1_ASAP7_75t_R _07860_ (.A(net3222),
    .B(_02126_),
    .Y(_02127_));
 OAI21x1_ASAP7_75t_R _07861_ (.A1(_02119_),
    .A2(_02126_),
    .B(_02093_),
    .Y(_02128_));
 OAI21x1_ASAP7_75t_R _07862_ (.A1(_02127_),
    .A2(_02128_),
    .B(net4163),
    .Y(_02129_));
 INVx1_ASAP7_75t_R _07863_ (.A(_02108_),
    .Y(_02130_));
 NAND2x1_ASAP7_75t_R _07864_ (.A(net3192),
    .B(net3181),
    .Y(_02131_));
 INVx1_ASAP7_75t_R _07865_ (.A(net3170),
    .Y(_02132_));
 OAI21x1_ASAP7_75t_R _07866_ (.A1(_02114_),
    .A2(_02102_),
    .B(_02078_),
    .Y(_02133_));
 XOR2x2_ASAP7_75t_R _07867_ (.A(net3144),
    .B(net4160),
    .Y(_02134_));
 NOR2x1_ASAP7_75t_R _07868_ (.A(_02132_),
    .B(_02134_),
    .Y(_02135_));
 AOI21x1_ASAP7_75t_R _07869_ (.A1(_02123_),
    .A2(net3184),
    .B(_02121_),
    .Y(_02136_));
 INVx1_ASAP7_75t_R _07870_ (.A(_02107_),
    .Y(_02137_));
 AOI21x1_ASAP7_75t_R _07871_ (.A1(_02129_),
    .A2(_02130_),
    .B(net3220),
    .Y(_02138_));
 NAND2x1_ASAP7_75t_R _07872_ (.A(_02137_),
    .B(_02138_),
    .Y(_02139_));
 OAI21x1_ASAP7_75t_R _07873_ (.A1(net3173),
    .A2(_02136_),
    .B(_02139_),
    .Y(_02140_));
 XOR2x2_ASAP7_75t_R _07874_ (.A(net3143),
    .B(net3182),
    .Y(_02141_));
 NAND2x1_ASAP7_75t_R _07875_ (.A(net3222),
    .B(net5440),
    .Y(_02142_));
 AO21x1_ASAP7_75t_R _07876_ (.A1(_02142_),
    .A2(_02093_),
    .B(net4163),
    .Y(_02143_));
 AOI21x1_ASAP7_75t_R _07877_ (.A1(net3220),
    .A2(_02143_),
    .B(_02099_),
    .Y(_02144_));
 INVx1_ASAP7_75t_R _07878_ (.A(net3169),
    .Y(_02145_));
 NOR2x1_ASAP7_75t_R _07879_ (.A(_02145_),
    .B(net3144),
    .Y(_02146_));
 OAI21x1_ASAP7_75t_R _07880_ (.A1(net3193),
    .A2(net3183),
    .B(_02137_),
    .Y(_02147_));
 XOR2x2_ASAP7_75t_R _07881_ (.A(net3169),
    .B(net3168),
    .Y(_02148_));
 AOI21x1_ASAP7_75t_R _07882_ (.A1(_02136_),
    .A2(_02139_),
    .B(net3173),
    .Y(_02149_));
 NOR2x1_ASAP7_75t_R _07883_ (.A(_02148_),
    .B(_02149_),
    .Y(_02150_));
 NOR2x1_ASAP7_75t_R _07884_ (.A(_02146_),
    .B(_02150_),
    .Y(_02151_));
 NAND2x1_ASAP7_75t_R _07885_ (.A(_02141_),
    .B(_02151_),
    .Y(_02152_));
 NOR2x1_ASAP7_75t_R _07886_ (.A(_02135_),
    .B(_02152_),
    .Y(_02153_));
 NAND2x1_ASAP7_75t_R _07887_ (.A(net4287),
    .B(net4376),
    .Y(_02154_));
 XOR2x2_ASAP7_75t_R _07888_ (.A(_02154_),
    .B(net4533),
    .Y(_02155_));
 INVx2_ASAP7_75t_R _07889_ (.A(_02155_),
    .Y(_02156_));
 OAI21x1_ASAP7_75t_R _07890_ (.A1(net3129),
    .A2(_02153_),
    .B(net4091),
    .Y(_02157_));
 XOR2x2_ASAP7_75t_R _07891_ (.A(net3172),
    .B(_02140_),
    .Y(_02158_));
 XNOR2x2_ASAP7_75t_R _07892_ (.A(_02144_),
    .B(_02147_),
    .Y(_02159_));
 NAND2x1_ASAP7_75t_R _07893_ (.A(_02159_),
    .B(_02133_),
    .Y(_02160_));
 NAND2x1_ASAP7_75t_R _07894_ (.A(net3169),
    .B(_02149_),
    .Y(_02161_));
 NAND2x1_ASAP7_75t_R _07895_ (.A(_02161_),
    .B(_02160_),
    .Y(_02162_));
 NOR2x2_ASAP7_75t_R _07896_ (.A(_02162_),
    .B(_02158_),
    .Y(_02163_));
 NOR3x1_ASAP7_75t_R _07897_ (.A(_02163_),
    .B(_02125_),
    .C(net4091),
    .Y(_02164_));
 INVx1_ASAP7_75t_R _07898_ (.A(_02164_),
    .Y(_02165_));
 OR2x2_ASAP7_75t_R _07899_ (.A(net4443),
    .B(net4342),
    .Y(_02166_));
 XOR2x2_ASAP7_75t_R _07900_ (.A(_02166_),
    .B(net4534),
    .Y(_02167_));
 INVx1_ASAP7_75t_R _07901_ (.A(_02167_),
    .Y(_02168_));
 NAND3x1_ASAP7_75t_R _07902_ (.A(_02157_),
    .B(_02165_),
    .C(_02168_),
    .Y(_02169_));
 INVx1_ASAP7_75t_R _07903_ (.A(_02125_),
    .Y(_02170_));
 XOR2x2_ASAP7_75t_R _07904_ (.A(_02133_),
    .B(net4092),
    .Y(_02171_));
 NAND2x1_ASAP7_75t_R _07905_ (.A(net3170),
    .B(_02171_),
    .Y(_02172_));
 NAND2x1_ASAP7_75t_R _07906_ (.A(_02172_),
    .B(_02163_),
    .Y(_02173_));
 AOI21x1_ASAP7_75t_R _07907_ (.A1(_02170_),
    .A2(_02173_),
    .B(net4158),
    .Y(_02174_));
 XOR2x2_ASAP7_75t_R _07908_ (.A(net3082),
    .B(net3128),
    .Y(_02175_));
 NAND3x1_ASAP7_75t_R _07909_ (.A(_02156_),
    .B(_02171_),
    .C(net3170),
    .Y(_02176_));
 OAI21x1_ASAP7_75t_R _07910_ (.A1(_02125_),
    .A2(net5397),
    .B(_02176_),
    .Y(_02177_));
 XOR2x2_ASAP7_75t_R _07911_ (.A(_02177_),
    .B(net3118),
    .Y(_02178_));
 NAND2x2_ASAP7_75t_R _07912_ (.A(_02171_),
    .B(_02156_),
    .Y(_02179_));
 XOR2x2_ASAP7_75t_R _07913_ (.A(_02131_),
    .B(net4160),
    .Y(_02180_));
 NOR2x1_ASAP7_75t_R _07914_ (.A(_02131_),
    .B(net3144),
    .Y(_02181_));
 AO21x1_ASAP7_75t_R _07915_ (.A1(net3144),
    .A2(_02180_),
    .B(_02181_),
    .Y(_02182_));
 AOI211x1_ASAP7_75t_R _07916_ (.A1(net5397),
    .A2(_02179_),
    .B(net3117),
    .C(net3130),
    .Y(_02183_));
 INVx1_ASAP7_75t_R _07917_ (.A(_02183_),
    .Y(_02184_));
 AOI21x1_ASAP7_75t_R _07918_ (.A1(net4091),
    .A2(_02135_),
    .B(_02152_),
    .Y(_02185_));
 XOR2x2_ASAP7_75t_R _07919_ (.A(_02182_),
    .B(_02179_),
    .Y(_02186_));
 OAI21x1_ASAP7_75t_R _07920_ (.A1(net3131),
    .A2(_02185_),
    .B(_02186_),
    .Y(_02187_));
 NAND2x2_ASAP7_75t_R _07921_ (.A(_02184_),
    .B(_02187_),
    .Y(_02188_));
 NOR2x2_ASAP7_75t_R _07922_ (.A(_02178_),
    .B(_02188_),
    .Y(_02189_));
 NAND2x1_ASAP7_75t_R _07923_ (.A(net3118),
    .B(_02176_),
    .Y(_02190_));
 OA21x2_ASAP7_75t_R _07924_ (.A1(_02190_),
    .A2(_02170_),
    .B(_02158_),
    .Y(_02191_));
 NOR2x2_ASAP7_75t_R _07925_ (.A(_02185_),
    .B(_02191_),
    .Y(_02192_));
 AOI21x1_ASAP7_75t_R _07926_ (.A1(_02175_),
    .A2(net3054),
    .B(net3080),
    .Y(_02193_));
 OAI21x1_ASAP7_75t_R _07927_ (.A1(net3073),
    .A2(_02193_),
    .B(net3072),
    .Y(_02194_));
 NOR3x1_ASAP7_75t_R _07928_ (.A(_02174_),
    .B(net4226),
    .C(net5382),
    .Y(_02195_));
 AND3x1_ASAP7_75t_R _07929_ (.A(_02192_),
    .B(net3127),
    .C(_02195_),
    .Y(_02196_));
 INVx1_ASAP7_75t_R _07930_ (.A(_02196_),
    .Y(_02197_));
 INVx1_ASAP7_75t_R _07931_ (.A(_02192_),
    .Y(_02198_));
 NOR2x1_ASAP7_75t_R _07932_ (.A(net3128),
    .B(_02169_),
    .Y(_02199_));
 OAI21x1_ASAP7_75t_R _07933_ (.A1(_02198_),
    .A2(_02199_),
    .B(net3071),
    .Y(_02200_));
 INVx2_ASAP7_75t_R _07934_ (.A(_02178_),
    .Y(_02201_));
 AOI21x1_ASAP7_75t_R _07935_ (.A1(net3127),
    .A2(_02195_),
    .B(_02188_),
    .Y(_02202_));
 OAI21x1_ASAP7_75t_R _07936_ (.A1(_02192_),
    .A2(_02201_),
    .B(_02202_),
    .Y(_02203_));
 NAND2x1_ASAP7_75t_R _07937_ (.A(_02203_),
    .B(_02200_),
    .Y(_02204_));
 AOI21x1_ASAP7_75t_R _07938_ (.A1(_02194_),
    .A2(_02197_),
    .B(_02204_),
    .Y(_02205_));
 AO21x1_ASAP7_75t_R _07939_ (.A1(_02176_),
    .A2(net5397),
    .B(net3131),
    .Y(_02206_));
 AOI21x1_ASAP7_75t_R _07940_ (.A1(net3107),
    .A2(_02206_),
    .B(net3096),
    .Y(_02207_));
 NAND2x1p5_ASAP7_75t_R _07941_ (.A(_02207_),
    .B(_02201_),
    .Y(_02208_));
 OAI21x1_ASAP7_75t_R _07942_ (.A1(_02208_),
    .A2(_02199_),
    .B(_02198_),
    .Y(_02209_));
 NAND2x1p5_ASAP7_75t_R _07943_ (.A(_02209_),
    .B(net4157),
    .Y(_02210_));
 NOR2x1_ASAP7_75t_R _07944_ (.A(_02164_),
    .B(_02174_),
    .Y(_02211_));
 NAND3x1_ASAP7_75t_R _07945_ (.A(_02211_),
    .B(net4156),
    .C(net3127),
    .Y(_02212_));
 AOI21x1_ASAP7_75t_R _07946_ (.A1(_02189_),
    .A2(_02212_),
    .B(_02192_),
    .Y(_02213_));
 NAND2x1_ASAP7_75t_R _07947_ (.A(net4226),
    .B(_02213_),
    .Y(_02214_));
 AND3x1_ASAP7_75t_R _07948_ (.A(net3084),
    .B(_01179_),
    .C(net3083),
    .Y(_02215_));
 NAND3x1_ASAP7_75t_R _07949_ (.A(_02210_),
    .B(_02214_),
    .C(_02215_),
    .Y(_02216_));
 NOR2x1_ASAP7_75t_R _07950_ (.A(_02208_),
    .B(_02199_),
    .Y(_02217_));
 AOI21x1_ASAP7_75t_R _07951_ (.A1(net3081),
    .A2(_02203_),
    .B(_02217_),
    .Y(_02218_));
 AOI21x1_ASAP7_75t_R _07952_ (.A1(_02205_),
    .A2(_02216_),
    .B(_02218_),
    .Y(_02219_));
 NAND2x1p5_ASAP7_75t_R _07953_ (.A(net4102),
    .B(_02219_),
    .Y(_02220_));
 INVx1_ASAP7_75t_R _07954_ (.A(_02175_),
    .Y(_02221_));
 AOI21x1_ASAP7_75t_R _07955_ (.A1(net3070),
    .A2(_02209_),
    .B(_02221_),
    .Y(_02222_));
 INVx1_ASAP7_75t_R _07956_ (.A(_02204_),
    .Y(_02223_));
 OAI21x1_ASAP7_75t_R _07957_ (.A1(net3053),
    .A2(_02222_),
    .B(_02223_),
    .Y(_02224_));
 INVx1_ASAP7_75t_R _07958_ (.A(_02215_),
    .Y(_02225_));
 XOR2x2_ASAP7_75t_R _07959_ (.A(net4157),
    .B(_02213_),
    .Y(_02226_));
 NOR2x2_ASAP7_75t_R _07960_ (.A(_02225_),
    .B(_02226_),
    .Y(_02227_));
 INVx1_ASAP7_75t_R _07961_ (.A(_02218_),
    .Y(_02228_));
 OAI21x1_ASAP7_75t_R _07962_ (.A1(_02224_),
    .A2(_02227_),
    .B(_02228_),
    .Y(_02229_));
 NAND2x2_ASAP7_75t_R _07963_ (.A(net5373),
    .B(net4177),
    .Y(_02230_));
 NAND2x1_ASAP7_75t_R _07964_ (.A(net2996),
    .B(net2983),
    .Y(_02231_));
 INVx1_ASAP7_75t_R _07965_ (.A(_02231_),
    .Y(_02232_));
 NOR2x1_ASAP7_75t_R _07966_ (.A(net4177),
    .B(net3026),
    .Y(_02233_));
 INVx1_ASAP7_75t_R _07967_ (.A(_02233_),
    .Y(_02234_));
 INVx1_ASAP7_75t_R _07968_ (.A(net3069),
    .Y(_02235_));
 NOR2x1_ASAP7_75t_R _07969_ (.A(net3073),
    .B(net3040),
    .Y(_02236_));
 AO21x1_ASAP7_75t_R _07970_ (.A1(net3029),
    .A2(_02235_),
    .B(_02236_),
    .Y(_02237_));
 OAI21x1_ASAP7_75t_R _07971_ (.A1(_02234_),
    .A2(_02219_),
    .B(_02237_),
    .Y(_02238_));
 NAND3x1_ASAP7_75t_R _07972_ (.A(net5373),
    .B(net3069),
    .C(_02233_),
    .Y(_02239_));
 NOR2x1_ASAP7_75t_R _07973_ (.A(_02196_),
    .B(_02222_),
    .Y(_02240_));
 NOR2x1_ASAP7_75t_R _07974_ (.A(_02240_),
    .B(_02227_),
    .Y(_02241_));
 INVx1_ASAP7_75t_R _07975_ (.A(_02240_),
    .Y(_02242_));
 AOI21x1_ASAP7_75t_R _07976_ (.A1(net3028),
    .A2(net3015),
    .B(_02242_),
    .Y(_02243_));
 AOI21x1_ASAP7_75t_R _07977_ (.A1(_02241_),
    .A2(_02229_),
    .B(_02243_),
    .Y(_02244_));
 INVx1_ASAP7_75t_R _07978_ (.A(_02244_),
    .Y(_02245_));
 AOI21x1_ASAP7_75t_R _07979_ (.A1(_02238_),
    .A2(_02239_),
    .B(_02245_),
    .Y(_02246_));
 AND2x2_ASAP7_75t_R _07980_ (.A(net4287),
    .B(net4479),
    .Y(_02247_));
 XNOR2x2_ASAP7_75t_R _07981_ (.A(net4538),
    .B(_02247_),
    .Y(_02248_));
 INVx1_ASAP7_75t_R _07982_ (.A(_02248_),
    .Y(_02249_));
 AOI21x1_ASAP7_75t_R _07983_ (.A1(_02220_),
    .A2(_02230_),
    .B(net3027),
    .Y(_02250_));
 NAND2x2_ASAP7_75t_R _07984_ (.A(_02250_),
    .B(_02249_),
    .Y(_02251_));
 NAND2x1_ASAP7_75t_R _07985_ (.A(_02241_),
    .B(net5373),
    .Y(_02252_));
 NAND2x1_ASAP7_75t_R _07986_ (.A(net3016),
    .B(net3015),
    .Y(_02253_));
 INVx1_ASAP7_75t_R _07987_ (.A(_02253_),
    .Y(_02254_));
 AOI21x1_ASAP7_75t_R _07988_ (.A1(net3030),
    .A2(_02252_),
    .B(_02254_),
    .Y(_02255_));
 AOI21x1_ASAP7_75t_R _07989_ (.A1(_02246_),
    .A2(_02251_),
    .B(_02255_),
    .Y(_02256_));
 XOR2x2_ASAP7_75t_R _07990_ (.A(_02256_),
    .B(net4090),
    .Y(_02257_));
 NOR2x1_ASAP7_75t_R _07991_ (.A(net2955),
    .B(_02257_),
    .Y(_02258_));
 AO21x1_ASAP7_75t_R _07992_ (.A1(net2983),
    .A2(net2996),
    .B(net4155),
    .Y(_02259_));
 NOR2x1_ASAP7_75t_R _07993_ (.A(net4177),
    .B(net3007),
    .Y(_02260_));
 XOR2x2_ASAP7_75t_R _07994_ (.A(_02260_),
    .B(net3027),
    .Y(_02261_));
 AOI21x1_ASAP7_75t_R _07995_ (.A1(_02261_),
    .A2(net5453),
    .B(net5421),
    .Y(_02262_));
 OAI21x1_ASAP7_75t_R _07996_ (.A1(_02259_),
    .A2(_02262_),
    .B(net2981),
    .Y(_02263_));
 INVx1_ASAP7_75t_R _07997_ (.A(_02263_),
    .Y(_02264_));
 NOR2x1_ASAP7_75t_R _07998_ (.A(net4102),
    .B(net3007),
    .Y(_02265_));
 NOR2x1_ASAP7_75t_R _07999_ (.A(net4177),
    .B(net5374),
    .Y(_02266_));
 INVx1_ASAP7_75t_R _08000_ (.A(net3027),
    .Y(_02267_));
 OAI21x1_ASAP7_75t_R _08001_ (.A1(_02265_),
    .A2(_02266_),
    .B(_02267_),
    .Y(_02268_));
 NOR2x1_ASAP7_75t_R _08002_ (.A(net4155),
    .B(_02268_),
    .Y(_02269_));
 INVx1_ASAP7_75t_R _08003_ (.A(_02238_),
    .Y(_02270_));
 NOR3x1_ASAP7_75t_R _08004_ (.A(_02219_),
    .B(net3052),
    .C(_02234_),
    .Y(_02271_));
 OAI21x1_ASAP7_75t_R _08005_ (.A1(_02270_),
    .A2(_02271_),
    .B(net2982),
    .Y(_02272_));
 INVx2_ASAP7_75t_R _08006_ (.A(_02255_),
    .Y(_02273_));
 OAI21x1_ASAP7_75t_R _08007_ (.A1(_02272_),
    .A2(_02269_),
    .B(_02273_),
    .Y(_02274_));
 NAND2x1_ASAP7_75t_R _08008_ (.A(_02274_),
    .B(_02269_),
    .Y(_02275_));
 INVx1_ASAP7_75t_R _08009_ (.A(_02275_),
    .Y(_02276_));
 OAI21x1_ASAP7_75t_R _08010_ (.A1(_02246_),
    .A2(_02255_),
    .B(_02251_),
    .Y(_02277_));
 NOR2x1_ASAP7_75t_R _08011_ (.A(_02270_),
    .B(_02271_),
    .Y(_02278_));
 XOR2x2_ASAP7_75t_R _08012_ (.A(net2969),
    .B(_02277_),
    .Y(_02279_));
 OAI21x1_ASAP7_75t_R _08013_ (.A1(_02264_),
    .A2(_02276_),
    .B(_02279_),
    .Y(_02280_));
 NAND2x1_ASAP7_75t_R _08014_ (.A(net2954),
    .B(net2953),
    .Y(_02281_));
 INVx1_ASAP7_75t_R _08015_ (.A(_02281_),
    .Y(_02282_));
 INVx1_ASAP7_75t_R _08016_ (.A(_02278_),
    .Y(_02283_));
 NAND2x1_ASAP7_75t_R _08017_ (.A(_02283_),
    .B(net2953),
    .Y(_02284_));
 OA21x2_ASAP7_75t_R _08018_ (.A1(_02284_),
    .A2(_02273_),
    .B(net2971),
    .Y(_02285_));
 NOR2x2_ASAP7_75t_R _08019_ (.A(_02282_),
    .B(_02285_),
    .Y(_02286_));
 INVx3_ASAP7_75t_R _08020_ (.A(_02286_),
    .Y(_02287_));
 OAI21x1_ASAP7_75t_R _08021_ (.A1(_02258_),
    .A2(_02280_),
    .B(_02287_),
    .Y(_02288_));
 NAND2x2_ASAP7_75t_R _08022_ (.A(_02288_),
    .B(net4103),
    .Y(_02289_));
 NAND2x1_ASAP7_75t_R _08023_ (.A(_02256_),
    .B(net4155),
    .Y(_02290_));
 NOR2x1_ASAP7_75t_R _08024_ (.A(net5451),
    .B(_02272_),
    .Y(_02291_));
 OAI21x1_ASAP7_75t_R _08025_ (.A1(net2970),
    .A2(_02291_),
    .B(net4090),
    .Y(_02292_));
 NAND3x1_ASAP7_75t_R _08026_ (.A(_02292_),
    .B(_02290_),
    .C(_01163_),
    .Y(_02293_));
 INVx1_ASAP7_75t_R _08027_ (.A(net2915),
    .Y(_02294_));
 XOR2x2_ASAP7_75t_R _08028_ (.A(_02231_),
    .B(net4090),
    .Y(_02295_));
 NAND2x1_ASAP7_75t_R _08029_ (.A(_02232_),
    .B(_02256_),
    .Y(_02296_));
 OAI21x1_ASAP7_75t_R _08030_ (.A1(_02295_),
    .A2(net2935),
    .B(_02296_),
    .Y(_02297_));
 NOR2x1_ASAP7_75t_R _08031_ (.A(_02293_),
    .B(_02297_),
    .Y(_02298_));
 OAI21x1_ASAP7_75t_R _08032_ (.A1(_02298_),
    .A2(net2892),
    .B(_02287_),
    .Y(_02299_));
 AOI22x1_ASAP7_75t_R _08033_ (.A1(net2926),
    .A2(_02289_),
    .B1(_02294_),
    .B2(_02299_),
    .Y(_02300_));
 XOR2x2_ASAP7_75t_R _08034_ (.A(net4155),
    .B(_02256_),
    .Y(_02301_));
 NAND2x1_ASAP7_75t_R _08035_ (.A(net2972),
    .B(_02301_),
    .Y(_02302_));
 AOI211x1_ASAP7_75t_R _08036_ (.A1(_02272_),
    .A2(_02273_),
    .B(net2952),
    .C(_02283_),
    .Y(_02303_));
 INVx1_ASAP7_75t_R _08037_ (.A(_02303_),
    .Y(_02304_));
 NAND2x1_ASAP7_75t_R _08038_ (.A(net2951),
    .B(net5448),
    .Y(_02305_));
 AOI22x1_ASAP7_75t_R _08039_ (.A1(_02263_),
    .A2(net5445),
    .B1(_02304_),
    .B2(_02305_),
    .Y(_02306_));
 NAND2x1_ASAP7_75t_R _08040_ (.A(_02302_),
    .B(_02306_),
    .Y(_02307_));
 AOI21x1_ASAP7_75t_R _08041_ (.A1(net2890),
    .A2(_02307_),
    .B(net4178),
    .Y(_02308_));
 NAND2x1_ASAP7_75t_R _08042_ (.A(net4582),
    .B(net4287),
    .Y(_02309_));
 XNOR2x2_ASAP7_75t_R _08043_ (.A(net4597),
    .B(_02309_),
    .Y(_02310_));
 INVx1_ASAP7_75t_R _08044_ (.A(_02310_),
    .Y(_02311_));
 NOR3x1_ASAP7_75t_R _08045_ (.A(net2913),
    .B(net4103),
    .C(net2916),
    .Y(_02312_));
 NOR3x2_ASAP7_75t_R _08046_ (.B(_02311_),
    .C(_02308_),
    .Y(_02313_),
    .A(_02312_));
 XOR2x2_ASAP7_75t_R _08047_ (.A(_02300_),
    .B(_02313_),
    .Y(_02314_));
 NAND2x1_ASAP7_75t_R _08048_ (.A(net5446),
    .B(net2925),
    .Y(_02315_));
 NAND3x2_ASAP7_75t_R _08049_ (.B(net4103),
    .C(net2972),
    .Y(_02316_),
    .A(_02301_));
 NAND2x1_ASAP7_75t_R _08050_ (.A(_02315_),
    .B(_02316_),
    .Y(_02317_));
 AOI21x1_ASAP7_75t_R _08051_ (.A1(net2912),
    .A2(_02316_),
    .B(net2916),
    .Y(_02318_));
 INVx1_ASAP7_75t_R _08052_ (.A(_02315_),
    .Y(_02319_));
 OAI21x1_ASAP7_75t_R _08053_ (.A1(net2891),
    .A2(net2889),
    .B(_02319_),
    .Y(_02320_));
 OAI21x1_ASAP7_75t_R _08054_ (.A1(net2888),
    .A2(_02318_),
    .B(_02320_),
    .Y(_02321_));
 XOR2x2_ASAP7_75t_R _08055_ (.A(_02293_),
    .B(_02297_),
    .Y(_02322_));
 INVx1_ASAP7_75t_R _08056_ (.A(_02322_),
    .Y(_02323_));
 INVx1_ASAP7_75t_R _08057_ (.A(net2914),
    .Y(_02324_));
 NOR3x1_ASAP7_75t_R _08058_ (.A(net2912),
    .B(net2916),
    .C(_02324_),
    .Y(_02325_));
 AOI21x1_ASAP7_75t_R _08059_ (.A1(_02323_),
    .A2(_02299_),
    .B(_02325_),
    .Y(_02326_));
 NOR2x1p5_ASAP7_75t_R _08060_ (.A(_02321_),
    .B(_02326_),
    .Y(_02327_));
 NAND2x1_ASAP7_75t_R _08061_ (.A(_02313_),
    .B(_02300_),
    .Y(_02328_));
 NAND2x1_ASAP7_75t_R _08062_ (.A(net2912),
    .B(net2910),
    .Y(_02329_));
 INVx1_ASAP7_75t_R _08063_ (.A(net2924),
    .Y(_02330_));
 OAI21x1_ASAP7_75t_R _08064_ (.A1(net2891),
    .A2(_02317_),
    .B(_02330_),
    .Y(_02331_));
 NAND2x2_ASAP7_75t_R _08065_ (.A(_02329_),
    .B(_02331_),
    .Y(_02332_));
 INVx1_ASAP7_75t_R _08066_ (.A(_02332_),
    .Y(_02333_));
 AOI21x1_ASAP7_75t_R _08067_ (.A1(net5769),
    .A2(_02328_),
    .B(_02333_),
    .Y(_02334_));
 NAND3x1_ASAP7_75t_R _08068_ (.A(net2892),
    .B(_02287_),
    .C(net2914),
    .Y(_02335_));
 OAI21x1_ASAP7_75t_R _08069_ (.A1(_02318_),
    .A2(_02322_),
    .B(_02335_),
    .Y(_02336_));
 NOR2x1_ASAP7_75t_R _08070_ (.A(_02319_),
    .B(_02298_),
    .Y(_02337_));
 AOI21x1_ASAP7_75t_R _08071_ (.A1(net2916),
    .A2(net2910),
    .B(net2911),
    .Y(_02338_));
 AOI21x1_ASAP7_75t_R _08072_ (.A1(_02337_),
    .A2(_02299_),
    .B(_02338_),
    .Y(_02339_));
 NAND2x2_ASAP7_75t_R _08073_ (.A(_02336_),
    .B(_02339_),
    .Y(_02340_));
 OAI22x1_ASAP7_75t_R _08074_ (.A1(net2877),
    .A2(net2923),
    .B1(net2915),
    .B2(net2887),
    .Y(_02341_));
 NAND3x1_ASAP7_75t_R _08075_ (.A(_02340_),
    .B(_02341_),
    .C(_02332_),
    .Y(_02342_));
 OAI21x1_ASAP7_75t_R _08076_ (.A1(_02314_),
    .A2(_02334_),
    .B(_02342_),
    .Y(_02343_));
 AOI22x1_ASAP7_75t_R _08077_ (.A1(_02340_),
    .A2(_02332_),
    .B1(net2847),
    .B2(_02313_),
    .Y(_02344_));
 XOR2x2_ASAP7_75t_R _08078_ (.A(_02344_),
    .B(net2861),
    .Y(_02345_));
 NOR2x1_ASAP7_75t_R _08079_ (.A(net5877),
    .B(_02345_),
    .Y(_02346_));
 AOI21x1_ASAP7_75t_R _08080_ (.A1(net2847),
    .A2(_02313_),
    .B(net5759),
    .Y(_02347_));
 NAND3x1_ASAP7_75t_R _08081_ (.A(net2893),
    .B(_02287_),
    .C(net4178),
    .Y(_02348_));
 NAND3x1_ASAP7_75t_R _08082_ (.A(net2923),
    .B(_02289_),
    .C(_02348_),
    .Y(_02349_));
 NOR2x1_ASAP7_75t_R _08083_ (.A(net4089),
    .B(_02349_),
    .Y(_02350_));
 OAI21x1_ASAP7_75t_R _08084_ (.A1(_02350_),
    .A2(_02340_),
    .B(_02332_),
    .Y(_02351_));
 NOR2x1_ASAP7_75t_R _08085_ (.A(_02312_),
    .B(net2877),
    .Y(_02352_));
 NAND2x1_ASAP7_75t_R _08086_ (.A(net4089),
    .B(_02352_),
    .Y(_02353_));
 NAND2x1_ASAP7_75t_R _08087_ (.A(net2861),
    .B(net5398),
    .Y(_02354_));
 NAND2x1_ASAP7_75t_R _08088_ (.A(net2861),
    .B(net2845),
    .Y(_02355_));
 OAI21x1_ASAP7_75t_R _08089_ (.A1(_02353_),
    .A2(_02354_),
    .B(_02355_),
    .Y(_02356_));
 AOI21x1_ASAP7_75t_R _08090_ (.A1(_02351_),
    .A2(_02356_),
    .B(net2860),
    .Y(_02357_));
 NOR2x1_ASAP7_75t_R _08091_ (.A(net2831),
    .B(_02357_),
    .Y(_02358_));
 OAI21x1_ASAP7_75t_R _08092_ (.A1(net4089),
    .A2(_02349_),
    .B(_02327_),
    .Y(_02359_));
 NAND3x1_ASAP7_75t_R _08093_ (.A(net2862),
    .B(net4089),
    .C(_02359_),
    .Y(_02360_));
 OAI21x1_ASAP7_75t_R _08094_ (.A1(net2846),
    .A2(_02347_),
    .B(net4154),
    .Y(_02361_));
 NAND2x1_ASAP7_75t_R _08095_ (.A(net4701),
    .B(net4287),
    .Y(_02362_));
 XOR2x2_ASAP7_75t_R _08096_ (.A(_02362_),
    .B(net4711),
    .Y(_02363_));
 INVx1_ASAP7_75t_R _08097_ (.A(_00466_),
    .Y(_02364_));
 NOR2x1_ASAP7_75t_R _08098_ (.A(net4598),
    .B(net4342),
    .Y(_02365_));
 XOR2x2_ASAP7_75t_R _08099_ (.A(_02365_),
    .B(net4596),
    .Y(_02366_));
 AND3x1_ASAP7_75t_R _08100_ (.A(_02363_),
    .B(_02364_),
    .C(_02366_),
    .Y(_02367_));
 AND3x1_ASAP7_75t_R _08101_ (.A(net2864),
    .B(_02367_),
    .C(net2876),
    .Y(_02368_));
 NAND3x1_ASAP7_75t_R _08102_ (.A(_02360_),
    .B(_02361_),
    .C(_02368_),
    .Y(_02369_));
 NOR2x1_ASAP7_75t_R _08103_ (.A(_02358_),
    .B(_02369_),
    .Y(_02370_));
 AOI21x1_ASAP7_75t_R _08104_ (.A1(_02346_),
    .A2(_02370_),
    .B(net4342),
    .Y(_02371_));
 BUFx3_ASAP7_75t_R place3021 (.A(_05157_),
    .Y(net3021));
 XOR2x2_ASAP7_75t_R _08106_ (.A(net2767),
    .B(net5114),
    .Y(_02373_));
 INVx1_ASAP7_75t_R _08107_ (.A(_02357_),
    .Y(_02374_));
 AO21x1_ASAP7_75t_R _08108_ (.A1(net2830),
    .A2(_02374_),
    .B(_02345_),
    .Y(_02375_));
 NOR2x1_ASAP7_75t_R _08109_ (.A(net4154),
    .B(_02351_),
    .Y(_02376_));
 AOI21x1_ASAP7_75t_R _08110_ (.A1(_02359_),
    .A2(net2862),
    .B(net4089),
    .Y(_02377_));
 AND3x1_ASAP7_75t_R _08111_ (.A(_02363_),
    .B(net5143),
    .C(_00465_),
    .Y(_02378_));
 AND2x2_ASAP7_75t_R _08112_ (.A(_02378_),
    .B(net4225),
    .Y(_02379_));
 INVx1_ASAP7_75t_R _08113_ (.A(_02379_),
    .Y(_02380_));
 NOR3x1_ASAP7_75t_R _08114_ (.A(_02380_),
    .B(_02377_),
    .C(_02376_),
    .Y(_02381_));
 OAI21x1_ASAP7_75t_R _08115_ (.A1(net4089),
    .A2(_02334_),
    .B(net2859),
    .Y(_02382_));
 INVx1_ASAP7_75t_R _08116_ (.A(net2859),
    .Y(_02383_));
 NAND2x1_ASAP7_75t_R _08117_ (.A(_02383_),
    .B(_02377_),
    .Y(_02384_));
 AOI21x1_ASAP7_75t_R _08118_ (.A1(_02382_),
    .A2(_02384_),
    .B(_02343_),
    .Y(_02385_));
 NAND2x1_ASAP7_75t_R _08119_ (.A(_02381_),
    .B(_02385_),
    .Y(_02386_));
 OAI21x1_ASAP7_75t_R _08120_ (.A1(_02386_),
    .A2(_02375_),
    .B(net4287),
    .Y(_02387_));
 BUFx3_ASAP7_75t_R place3020 (.A(_05190_),
    .Y(net3020));
 INVx1_ASAP7_75t_R _08122_ (.A(_00032_),
    .Y(_02389_));
 XOR2x2_ASAP7_75t_R _08123_ (.A(net5394),
    .B(net5015),
    .Y(_02390_));
 NAND2x1_ASAP7_75t_R _08124_ (.A(_02373_),
    .B(_02390_),
    .Y(_02391_));
 INVx1_ASAP7_75t_R _08125_ (.A(net5083),
    .Y(_02392_));
 XOR2x1_ASAP7_75t_R _08126_ (.A(net5014),
    .Y(_02393_),
    .B(net2765));
 NAND2x1_ASAP7_75t_R _08127_ (.A(net2830),
    .B(net2794),
    .Y(_02394_));
 INVx1_ASAP7_75t_R _08128_ (.A(net2844),
    .Y(_02395_));
 NAND2x1_ASAP7_75t_R _08129_ (.A(net2819),
    .B(net2820),
    .Y(_02396_));
 NOR2x1_ASAP7_75t_R _08130_ (.A(_02395_),
    .B(_02396_),
    .Y(_02397_));
 AOI21x1_ASAP7_75t_R _08131_ (.A1(net2796),
    .A2(_02397_),
    .B(net4342),
    .Y(_02398_));
 NAND2x1_ASAP7_75t_R _08132_ (.A(_02394_),
    .B(_02398_),
    .Y(_02399_));
 INVx1_ASAP7_75t_R _08133_ (.A(_02314_),
    .Y(_02400_));
 INVx1_ASAP7_75t_R _08134_ (.A(net2833),
    .Y(_02401_));
 AOI21x1_ASAP7_75t_R _08135_ (.A1(net2821),
    .A2(_02400_),
    .B(_02401_),
    .Y(_02402_));
 XOR2x2_ASAP7_75t_R _08136_ (.A(net2832),
    .B(net2863),
    .Y(_02403_));
 NAND2x1_ASAP7_75t_R _08137_ (.A(_02402_),
    .B(_02403_),
    .Y(_02404_));
 OAI21x1_ASAP7_75t_R _08138_ (.A1(net2809),
    .A2(_02404_),
    .B(net4287),
    .Y(_02405_));
 NAND2x1_ASAP7_75t_R _08139_ (.A(net2795),
    .B(_02405_),
    .Y(_02406_));
 INVx2_ASAP7_75t_R _08140_ (.A(_00029_),
    .Y(_02407_));
 NAND3x1_ASAP7_75t_R _08141_ (.A(_02399_),
    .B(_02406_),
    .C(net5013),
    .Y(_02408_));
 NOR2x1_ASAP7_75t_R _08142_ (.A(net2795),
    .B(_02405_),
    .Y(_02409_));
 INVx1_ASAP7_75t_R _08143_ (.A(_02406_),
    .Y(_02410_));
 OAI21x1_ASAP7_75t_R _08144_ (.A1(_02409_),
    .A2(_02410_),
    .B(net5084),
    .Y(_02411_));
 NAND3x1_ASAP7_75t_R _08145_ (.A(_02411_),
    .B(_02408_),
    .C(_02393_),
    .Y(_02412_));
 NOR2x1_ASAP7_75t_R _08146_ (.A(_02391_),
    .B(_02412_),
    .Y(_02413_));
 XOR2x2_ASAP7_75t_R _08147_ (.A(net2810),
    .B(net5086),
    .Y(_02414_));
 NAND2x1_ASAP7_75t_R _08148_ (.A(net4287),
    .B(net2809),
    .Y(_02415_));
 XNOR2x2_ASAP7_75t_R _08149_ (.A(_02414_),
    .B(_02415_),
    .Y(_02416_));
 AO21x1_ASAP7_75t_R _08150_ (.A1(_02385_),
    .A2(net2793),
    .B(net4342),
    .Y(_02417_));
 XOR2x2_ASAP7_75t_R _08151_ (.A(_02403_),
    .B(net5085),
    .Y(_02418_));
 XOR2x2_ASAP7_75t_R _08152_ (.A(_02417_),
    .B(_02418_),
    .Y(_02419_));
 NAND2x1_ASAP7_75t_R _08153_ (.A(_02416_),
    .B(_02419_),
    .Y(_02420_));
 NOR2x1_ASAP7_75t_R _08154_ (.A(net4342),
    .B(net4022),
    .Y(_02421_));
 BUFx3_ASAP7_75t_R place3018 (.A(_06262_),
    .Y(net3018));
 XOR2x2_ASAP7_75t_R _08156_ (.A(_02421_),
    .B(net5087),
    .Y(_02423_));
 XOR2x2_ASAP7_75t_R _08157_ (.A(net2806),
    .B(_02423_),
    .Y(_02424_));
 NAND2x1_ASAP7_75t_R _08158_ (.A(net2808),
    .B(net2807),
    .Y(_02425_));
 INVx1_ASAP7_75t_R _08159_ (.A(_00026_),
    .Y(_02426_));
 XOR2x2_ASAP7_75t_R _08160_ (.A(_02425_),
    .B(net5012),
    .Y(_02427_));
 NOR2x1_ASAP7_75t_R _08161_ (.A(net4342),
    .B(net2793),
    .Y(_02428_));
 XOR2x2_ASAP7_75t_R _08162_ (.A(_02427_),
    .B(_02428_),
    .Y(_02429_));
 NAND2x1_ASAP7_75t_R _08163_ (.A(_02424_),
    .B(_02429_),
    .Y(_02430_));
 NOR2x1_ASAP7_75t_R _08164_ (.A(net4342),
    .B(net4088),
    .Y(_02431_));
 XOR2x2_ASAP7_75t_R _08165_ (.A(net4225),
    .B(net5089),
    .Y(_02432_));
 XOR2x2_ASAP7_75t_R _08166_ (.A(_02431_),
    .B(_02432_),
    .Y(_02433_));
 AO21x1_ASAP7_75t_R _08167_ (.A1(_00467_),
    .A2(net4287),
    .B(net4236),
    .Y(_02434_));
 XNOR2x2_ASAP7_75t_R _08168_ (.A(net5143),
    .B(net5635),
    .Y(_02435_));
 OAI21x1_ASAP7_75t_R _08169_ (.A1(net5020),
    .A2(_02434_),
    .B(_02435_),
    .Y(_02436_));
 AO21x1_ASAP7_75t_R _08170_ (.A1(net5020),
    .A2(_02434_),
    .B(_02436_),
    .Y(_02437_));
 NOR2x1_ASAP7_75t_R _08171_ (.A(net4046),
    .B(net4342),
    .Y(_02438_));
 XOR2x2_ASAP7_75t_R _08172_ (.A(_02438_),
    .B(net5092),
    .Y(_02439_));
 XNOR2x2_ASAP7_75t_R _08173_ (.A(_02439_),
    .B(net4153),
    .Y(_02440_));
 INVx1_ASAP7_75t_R _08174_ (.A(_02440_),
    .Y(_02441_));
 OR3x1_ASAP7_75t_R _08175_ (.A(_02433_),
    .B(_02437_),
    .C(_02441_),
    .Y(_02442_));
 NOR3x1_ASAP7_75t_R _08176_ (.A(_02420_),
    .B(_02430_),
    .C(_02442_),
    .Y(_02443_));
 XOR2x2_ASAP7_75t_R _08177_ (.A(net2767),
    .B(net5110),
    .Y(_02444_));
 INVx1_ASAP7_75t_R _08178_ (.A(_00036_),
    .Y(_02445_));
 XOR2x1_ASAP7_75t_R _08179_ (.A(net2766),
    .Y(_02446_),
    .B(net5011));
 NAND2x1_ASAP7_75t_R _08180_ (.A(_02444_),
    .B(_02446_),
    .Y(_02447_));
 XOR2x2_ASAP7_75t_R _08181_ (.A(net2767),
    .B(net5112),
    .Y(_02448_));
 INVx1_ASAP7_75t_R _08182_ (.A(_00034_),
    .Y(_02449_));
 XOR2x1_ASAP7_75t_R _08183_ (.A(net2766),
    .Y(_02450_),
    .B(net5009));
 NAND2x1_ASAP7_75t_R _08184_ (.A(_02448_),
    .B(_02450_),
    .Y(_02451_));
 NOR2x1_ASAP7_75t_R _08185_ (.A(_02451_),
    .B(_02447_),
    .Y(_02452_));
 NAND3x1_ASAP7_75t_R _08186_ (.A(_02452_),
    .B(_02443_),
    .C(_02413_),
    .Y(_02453_));
 INVx1_ASAP7_75t_R _08187_ (.A(net5096),
    .Y(_02454_));
 XOR2x2_ASAP7_75t_R _08188_ (.A(net2767),
    .B(net5008),
    .Y(_02455_));
 XOR2x2_ASAP7_75t_R _08189_ (.A(net2765),
    .B(net5095),
    .Y(_02456_));
 NOR2x1_ASAP7_75t_R _08190_ (.A(_02455_),
    .B(_02456_),
    .Y(_02457_));
 INVx1_ASAP7_75t_R _08191_ (.A(_00045_),
    .Y(_02458_));
 XOR2x2_ASAP7_75t_R _08192_ (.A(net2767),
    .B(net5007),
    .Y(_02459_));
 XOR2x2_ASAP7_75t_R _08193_ (.A(net2765),
    .B(net5098),
    .Y(_02460_));
 NOR2x1_ASAP7_75t_R _08194_ (.A(_02459_),
    .B(_02460_),
    .Y(_02461_));
 NAND2x1_ASAP7_75t_R _08195_ (.A(_02457_),
    .B(_02461_),
    .Y(_02462_));
 INVx1_ASAP7_75t_R _08196_ (.A(_00052_),
    .Y(_02463_));
 XOR2x2_ASAP7_75t_R _08197_ (.A(net2767),
    .B(net5006),
    .Y(_02464_));
 XOR2x2_ASAP7_75t_R _08198_ (.A(net2765),
    .B(net5090),
    .Y(_02465_));
 NOR2x1_ASAP7_75t_R _08199_ (.A(_02464_),
    .B(_02465_),
    .Y(_02466_));
 NAND2x1_ASAP7_75t_R _08200_ (.A(net5094),
    .B(net5394),
    .Y(_02467_));
 OR2x2_ASAP7_75t_R _08201_ (.A(net5094),
    .B(net5394),
    .Y(_02468_));
 INVx1_ASAP7_75t_R _08202_ (.A(_00050_),
    .Y(_02469_));
 XOR2x2_ASAP7_75t_R _08203_ (.A(net2767),
    .B(net5005),
    .Y(_02470_));
 AOI21x1_ASAP7_75t_R _08204_ (.A1(_02467_),
    .A2(_02468_),
    .B(_02470_),
    .Y(_02471_));
 NAND2x1_ASAP7_75t_R _08205_ (.A(_02466_),
    .B(_02471_),
    .Y(_02472_));
 NOR2x1_ASAP7_75t_R _08206_ (.A(_02472_),
    .B(_02462_),
    .Y(_02473_));
 XNOR2x2_ASAP7_75t_R _08207_ (.A(net5106),
    .B(net2767),
    .Y(_02474_));
 XOR2x2_ASAP7_75t_R _08208_ (.A(net2765),
    .B(net5105),
    .Y(_02475_));
 NOR2x1_ASAP7_75t_R _08209_ (.A(_02474_),
    .B(_02475_),
    .Y(_02476_));
 INVx1_ASAP7_75t_R _08210_ (.A(_00037_),
    .Y(_02477_));
 XOR2x2_ASAP7_75t_R _08211_ (.A(net2767),
    .B(net5004),
    .Y(_02478_));
 XOR2x1_ASAP7_75t_R _08212_ (.A(net5107),
    .Y(_02479_),
    .B(net2765));
 NOR2x1_ASAP7_75t_R _08213_ (.A(_02478_),
    .B(_02479_),
    .Y(_02480_));
 NAND2x1_ASAP7_75t_R _08214_ (.A(_02476_),
    .B(_02480_),
    .Y(_02481_));
 XNOR2x2_ASAP7_75t_R _08215_ (.A(net5103),
    .B(net2767),
    .Y(_02482_));
 XOR2x1_ASAP7_75t_R _08216_ (.A(net5394),
    .Y(_02483_),
    .B(net5102));
 NOR2x1_ASAP7_75t_R _08217_ (.A(_02482_),
    .B(_02483_),
    .Y(_02484_));
 OR2x2_ASAP7_75t_R _08218_ (.A(net5100),
    .B(net5394),
    .Y(_02485_));
 NAND2x1_ASAP7_75t_R _08219_ (.A(net5100),
    .B(net5394),
    .Y(_02486_));
 INVx1_ASAP7_75t_R _08220_ (.A(_00043_),
    .Y(_02487_));
 XOR2x2_ASAP7_75t_R _08221_ (.A(net2767),
    .B(net5003),
    .Y(_02488_));
 AOI21x1_ASAP7_75t_R _08222_ (.A1(_02485_),
    .A2(_02486_),
    .B(_02488_),
    .Y(_02489_));
 NAND2x1_ASAP7_75t_R _08223_ (.A(_02484_),
    .B(_02489_),
    .Y(_02490_));
 NOR2x1_ASAP7_75t_R _08224_ (.A(_02490_),
    .B(_02481_),
    .Y(_02491_));
 NAND2x1p5_ASAP7_75t_R _08225_ (.A(_02473_),
    .B(_02491_),
    .Y(_02492_));
 OA22x2_ASAP7_75t_R _08226_ (.A1(_01134_),
    .A2(_01143_),
    .B1(_02453_),
    .B2(net2725),
    .Y(_00023_));
 INVx1_ASAP7_75t_R _08227_ (.A(_00470_),
    .Y(\u_dct.k_ptr[0] ));
 INVx1_ASAP7_75t_R _08228_ (.A(_00471_),
    .Y(\u_dct.k_ptr[1] ));
 INVx1_ASAP7_75t_R _08229_ (.A(_00475_),
    .Y(\u_dct.n_ptr[0] ));
 INVx1_ASAP7_75t_R _08230_ (.A(_00476_),
    .Y(\u_dct.n_ptr[1] ));
 INVx1_ASAP7_75t_R _08231_ (.A(_00486_),
    .Y(_00487_));
 INVx1_ASAP7_75t_R _08232_ (.A(_00066_),
    .Y(\u_fft.sched[47] ));
 INVx1_ASAP7_75t_R _08233_ (.A(_00226_),
    .Y(\u_fft.sched[46] ));
 INVx1_ASAP7_75t_R _08234_ (.A(_00225_),
    .Y(\u_fft.sched[48] ));
 INVx1_ASAP7_75t_R _08235_ (.A(_00065_),
    .Y(\u_fft.sched[49] ));
 INVx1_ASAP7_75t_R _08236_ (.A(_00064_),
    .Y(\u_fft.sched[50] ));
 INVx1_ASAP7_75t_R _08237_ (.A(_00063_),
    .Y(\u_fft.sched[51] ));
 INVx1_ASAP7_75t_R _08238_ (.A(_00224_),
    .Y(\u_fft.sched[52] ));
 INVx1_ASAP7_75t_R _08239_ (.A(_00062_),
    .Y(\u_fft.sched[53] ));
 INVx1_ASAP7_75t_R _08240_ (.A(_00497_),
    .Y(_00338_));
 INVx1_ASAP7_75t_R _08241_ (.A(_00215_),
    .Y(\u_fft.sched[64] ));
 INVx1_ASAP7_75t_R _08242_ (.A(_00293_),
    .Y(\u_fft.power_ptr[0] ));
 INVx1_ASAP7_75t_R _08243_ (.A(_00292_),
    .Y(\u_fft.power_ptr[1] ));
 INVx1_ASAP7_75t_R _08244_ (.A(net5221),
    .Y(\u_hamming_window.frame_ptr[0] ));
 INVx1_ASAP7_75t_R _08245_ (.A(_00519_),
    .Y(\mel_ptr[1] ));
 INVx2_ASAP7_75t_R _08246_ (.A(_00518_),
    .Y(\mel_ptr[0] ));
 INVx1_ASAP7_75t_R _08247_ (.A(_00140_),
    .Y(\u_window_buffer.internal_read_ptr[30] ));
 INVx1_ASAP7_75t_R _08248_ (.A(_00141_),
    .Y(\u_window_buffer.internal_read_ptr[29] ));
 INVx1_ASAP7_75t_R _08249_ (.A(_00142_),
    .Y(\u_window_buffer.internal_read_ptr[28] ));
 INVx1_ASAP7_75t_R _08250_ (.A(_00143_),
    .Y(\u_window_buffer.internal_read_ptr[27] ));
 INVx2_ASAP7_75t_R _08251_ (.A(_00144_),
    .Y(\u_window_buffer.internal_read_ptr[26] ));
 INVx2_ASAP7_75t_R _08252_ (.A(_00145_),
    .Y(\u_window_buffer.internal_read_ptr[25] ));
 INVx2_ASAP7_75t_R _08253_ (.A(_00146_),
    .Y(\u_window_buffer.internal_read_ptr[24] ));
 INVx1_ASAP7_75t_R _08254_ (.A(_00147_),
    .Y(\u_window_buffer.internal_read_ptr[23] ));
 INVx2_ASAP7_75t_R _08255_ (.A(_00148_),
    .Y(\u_window_buffer.internal_read_ptr[22] ));
 INVx2_ASAP7_75t_R _08256_ (.A(_00149_),
    .Y(\u_window_buffer.internal_read_ptr[21] ));
 INVx2_ASAP7_75t_R _08257_ (.A(_00150_),
    .Y(\u_window_buffer.internal_read_ptr[20] ));
 INVx2_ASAP7_75t_R _08258_ (.A(_00151_),
    .Y(\u_window_buffer.internal_read_ptr[19] ));
 INVx2_ASAP7_75t_R _08259_ (.A(_00152_),
    .Y(\u_window_buffer.internal_read_ptr[18] ));
 INVx2_ASAP7_75t_R _08260_ (.A(_00153_),
    .Y(\u_window_buffer.internal_read_ptr[17] ));
 INVx2_ASAP7_75t_R _08261_ (.A(_00154_),
    .Y(\u_window_buffer.internal_read_ptr[16] ));
 INVx2_ASAP7_75t_R _08262_ (.A(_00155_),
    .Y(\u_window_buffer.internal_read_ptr[15] ));
 INVx2_ASAP7_75t_R _08263_ (.A(_00156_),
    .Y(\u_window_buffer.internal_read_ptr[14] ));
 INVx2_ASAP7_75t_R _08264_ (.A(_00157_),
    .Y(\u_window_buffer.internal_read_ptr[13] ));
 INVx2_ASAP7_75t_R _08265_ (.A(_00158_),
    .Y(\u_window_buffer.internal_read_ptr[12] ));
 INVx1_ASAP7_75t_R _08266_ (.A(_00159_),
    .Y(\u_window_buffer.internal_read_ptr[11] ));
 INVx3_ASAP7_75t_R _08267_ (.A(_00160_),
    .Y(\u_window_buffer.internal_read_ptr[10] ));
 INVx2_ASAP7_75t_R _08268_ (.A(_00134_),
    .Y(\u_window_buffer.internal_read_ptr[9] ));
 INVx1_ASAP7_75t_R _08269_ (.A(_00135_),
    .Y(\u_window_buffer.internal_read_ptr[8] ));
 INVx4_ASAP7_75t_R _08270_ (.A(_00136_),
    .Y(\u_window_buffer.internal_read_ptr[7] ));
 INVx2_ASAP7_75t_R _08271_ (.A(_00523_),
    .Y(\u_window_buffer.internal_read_ptr[1] ));
 INVx1_ASAP7_75t_R _08272_ (.A(net5177),
    .Y(_02493_));
 OR4x1_ASAP7_75t_R _08273_ (.A(net5178),
    .B(net5180),
    .C(net5181),
    .D(net5182),
    .Y(_02494_));
 AOI21x1_ASAP7_75t_R _08274_ (.A1(net5173),
    .A2(_00533_),
    .B(net5172),
    .Y(_02495_));
 AND3x4_ASAP7_75t_R _08275_ (.A(_02495_),
    .B(net4973),
    .C(net4974),
    .Y(_02496_));
 AND3x4_ASAP7_75t_R _08276_ (.A(_02496_),
    .B(net4976),
    .C(net4975),
    .Y(_02497_));
 NOR2x1_ASAP7_75t_R _08277_ (.A(net5193),
    .B(net5194),
    .Y(_02498_));
 AND3x1_ASAP7_75t_R _08278_ (.A(_02498_),
    .B(net4978),
    .C(net4977),
    .Y(_02499_));
 AND5x1_ASAP7_75t_R _08279_ (.A(net4984),
    .B(_02499_),
    .C(net4983),
    .D(net4982),
    .E(net4981),
    .Y(_02500_));
 NAND2x2_ASAP7_75t_R _08280_ (.A(net4639),
    .B(_02500_),
    .Y(_02501_));
 OR2x2_ASAP7_75t_R _08281_ (.A(net5188),
    .B(_02501_),
    .Y(_02502_));
 OR4x1_ASAP7_75t_R _08282_ (.A(net5183),
    .B(net5184),
    .C(net5185),
    .D(net5186),
    .Y(_02503_));
 OR3x1_ASAP7_75t_R _08283_ (.A(_02503_),
    .B(net5187),
    .C(_02502_),
    .Y(_02504_));
 NOR2x1_ASAP7_75t_R _08284_ (.A(_02504_),
    .B(_02494_),
    .Y(_02505_));
 NOR2x1p5_ASAP7_75t_R _08285_ (.A(_02493_),
    .B(_02505_),
    .Y(_02506_));
 AND2x4_ASAP7_75t_R _08286_ (.A(_02505_),
    .B(_02493_),
    .Y(_02507_));
 NOR2x1p5_ASAP7_75t_R _08287_ (.A(_02507_),
    .B(_02506_),
    .Y(_02508_));
 BUFx3_ASAP7_75t_R place3017 (.A(_06304_),
    .Y(net3017));
 BUFx3_ASAP7_75t_R place3016 (.A(_02205_),
    .Y(net3016));
 INVx2_ASAP7_75t_R _08290_ (.A(_00524_),
    .Y(\u_window_buffer.internal_read_ptr[2] ));
 NOR2x2_ASAP7_75t_R _08291_ (.A(net4968),
    .B(net4330),
    .Y(_02511_));
 AO21x1_ASAP7_75t_R _08292_ (.A1(_00526_),
    .A2(net4330),
    .B(_02511_),
    .Y(_00528_));
 INVx2_ASAP7_75t_R _08293_ (.A(_00058_),
    .Y(\u_window_buffer.internal_read_ptr[3] ));
 INVx1_ASAP7_75t_R _08294_ (.A(_00059_),
    .Y(\u_window_buffer.internal_read_ptr[4] ));
 INVx3_ASAP7_75t_R _08295_ (.A(_00138_),
    .Y(\u_window_buffer.internal_read_ptr[5] ));
 INVx2_ASAP7_75t_R _08296_ (.A(_00137_),
    .Y(\u_window_buffer.internal_read_ptr[6] ));
 INVx1_ASAP7_75t_R _08297_ (.A(net5171),
    .Y(\u_window_buffer.move_counter[0] ));
 INVx1_ASAP7_75t_R _08298_ (.A(_00081_),
    .Y(\u_window_buffer.read_ptr[30] ));
 INVx1_ASAP7_75t_R _08299_ (.A(_00083_),
    .Y(\u_window_buffer.read_ptr[29] ));
 INVx1_ASAP7_75t_R _08300_ (.A(_00084_),
    .Y(\u_window_buffer.read_ptr[28] ));
 INVx1_ASAP7_75t_R _08301_ (.A(_00085_),
    .Y(\u_window_buffer.read_ptr[27] ));
 INVx1_ASAP7_75t_R _08302_ (.A(_00086_),
    .Y(\u_window_buffer.read_ptr[26] ));
 INVx1_ASAP7_75t_R _08303_ (.A(_00087_),
    .Y(\u_window_buffer.read_ptr[25] ));
 INVx2_ASAP7_75t_R _08304_ (.A(_00088_),
    .Y(\u_window_buffer.read_ptr[24] ));
 INVx1_ASAP7_75t_R _08305_ (.A(_00089_),
    .Y(\u_window_buffer.read_ptr[23] ));
 INVx2_ASAP7_75t_R _08306_ (.A(_00090_),
    .Y(\u_window_buffer.read_ptr[22] ));
 INVx1_ASAP7_75t_R _08307_ (.A(_00091_),
    .Y(\u_window_buffer.read_ptr[21] ));
 INVx2_ASAP7_75t_R _08308_ (.A(_00092_),
    .Y(\u_window_buffer.read_ptr[20] ));
 INVx1_ASAP7_75t_R _08309_ (.A(_00094_),
    .Y(\u_window_buffer.read_ptr[19] ));
 INVx2_ASAP7_75t_R _08310_ (.A(_00095_),
    .Y(\u_window_buffer.read_ptr[18] ));
 INVx2_ASAP7_75t_R _08311_ (.A(_00096_),
    .Y(\u_window_buffer.read_ptr[17] ));
 INVx2_ASAP7_75t_R _08312_ (.A(_00097_),
    .Y(\u_window_buffer.read_ptr[16] ));
 INVx2_ASAP7_75t_R _08313_ (.A(_00098_),
    .Y(\u_window_buffer.read_ptr[15] ));
 INVx2_ASAP7_75t_R _08314_ (.A(_00099_),
    .Y(\u_window_buffer.read_ptr[14] ));
 INVx2_ASAP7_75t_R _08315_ (.A(_00100_),
    .Y(\u_window_buffer.read_ptr[13] ));
 INVx2_ASAP7_75t_R _08316_ (.A(_00101_),
    .Y(\u_window_buffer.read_ptr[12] ));
 INVx1_ASAP7_75t_R _08317_ (.A(_00102_),
    .Y(\u_window_buffer.read_ptr[11] ));
 INVx2_ASAP7_75t_R _08318_ (.A(_00103_),
    .Y(\u_window_buffer.read_ptr[10] ));
 INVx1_ASAP7_75t_R _08319_ (.A(_00073_),
    .Y(\u_window_buffer.read_ptr[9] ));
 INVx2_ASAP7_75t_R _08320_ (.A(_00074_),
    .Y(\u_window_buffer.read_ptr[8] ));
 INVx2_ASAP7_75t_R _08321_ (.A(_00075_),
    .Y(\u_window_buffer.read_ptr[7] ));
 INVx2_ASAP7_75t_R _08322_ (.A(_00076_),
    .Y(\u_window_buffer.read_ptr[6] ));
 INVx1_ASAP7_75t_R _08323_ (.A(_00077_),
    .Y(\u_window_buffer.read_ptr[5] ));
 INVx1_ASAP7_75t_R _08324_ (.A(_00078_),
    .Y(\u_window_buffer.read_ptr[4] ));
 INVx1_ASAP7_75t_R _08325_ (.A(_00079_),
    .Y(\u_window_buffer.read_ptr[3] ));
 INVx2_ASAP7_75t_R _08326_ (.A(_00082_),
    .Y(\u_window_buffer.read_ptr[2] ));
 INVx1_ASAP7_75t_R _08327_ (.A(_00093_),
    .Y(\u_window_buffer.read_ptr[1] ));
 BUFx3_ASAP7_75t_R place3019 (.A(_06262_),
    .Y(net3019));
 OR4x1_ASAP7_75t_R _08329_ (.A(_00951_),
    .B(_00177_),
    .C(_00326_),
    .D(_00328_),
    .Y(_02513_));
 NOR2x1_ASAP7_75t_R _08330_ (.A(net5360),
    .B(net4690),
    .Y(_00003_));
 INVx1_ASAP7_75t_R _08331_ (.A(_00936_),
    .Y(_02514_));
 BUFx3_ASAP7_75t_R place3015 (.A(_02216_),
    .Y(net3015));
 AND3x1_ASAP7_75t_R _08333_ (.A(_02514_),
    .B(net5362),
    .C(net5047),
    .Y(_00000_));
 INVx1_ASAP7_75t_R _08334_ (.A(_00941_),
    .Y(_02516_));
 AND3x1_ASAP7_75t_R _08335_ (.A(_02516_),
    .B(net5362),
    .C(net5045),
    .Y(_00001_));
 INVx1_ASAP7_75t_R _08336_ (.A(net5205),
    .Y(_02517_));
 AND3x1_ASAP7_75t_R _08337_ (.A(net4751),
    .B(net4934),
    .C(_00902_),
    .Y(_00004_));
 INVx1_ASAP7_75t_R _08338_ (.A(_00324_),
    .Y(_02518_));
 AND3x1_ASAP7_75t_R _08339_ (.A(net4933),
    .B(net5362),
    .C(net4746),
    .Y(_00002_));
 INVx1_ASAP7_75t_R _08340_ (.A(_00549_),
    .Y(\u_hamming_window.calc_pointer[1] ));
 INVx1_ASAP7_75t_R _08341_ (.A(_00548_),
    .Y(\u_hamming_window.calc_pointer[0] ));
 INVx1_ASAP7_75t_R _08342_ (.A(net5211),
    .Y(\u_mel.k[1] ));
 INVx1_ASAP7_75t_R _08343_ (.A(\u_mel.k_next[0] ),
    .Y(\u_mel.k[0] ));
 INVx1_ASAP7_75t_R _08344_ (.A(_00216_),
    .Y(\u_fft.sched[63] ));
 INVx1_ASAP7_75t_R _08345_ (.A(_00217_),
    .Y(\u_fft.sched[62] ));
 INVx1_ASAP7_75t_R _08346_ (.A(_00218_),
    .Y(\u_fft.sched[61] ));
 INVx1_ASAP7_75t_R _08347_ (.A(_00219_),
    .Y(\u_fft.sched[60] ));
 INVx1_ASAP7_75t_R _08348_ (.A(_00220_),
    .Y(\u_fft.sched[59] ));
 INVx1_ASAP7_75t_R _08349_ (.A(_00221_),
    .Y(\u_fft.sched[58] ));
 INVx1_ASAP7_75t_R _08350_ (.A(_00222_),
    .Y(\u_fft.sched[57] ));
 INVx1_ASAP7_75t_R _08351_ (.A(_00223_),
    .Y(\u_fft.sched[56] ));
 INVx1_ASAP7_75t_R _08352_ (.A(_00494_),
    .Y(\u_fft.sched[55] ));
 INVx1_ASAP7_75t_R _08353_ (.A(_00061_),
    .Y(\u_fft.sched[54] ));
 INVx1_ASAP7_75t_R _08354_ (.A(_00318_),
    .Y(net213));
 INVx1_ASAP7_75t_R _08355_ (.A(_00325_),
    .Y(\u_hamming_window.done ));
 AO21x1_ASAP7_75t_R _08356_ (.A1(_00046_),
    .A2(net5213),
    .B(_01008_),
    .Y(_02519_));
 INVx1_ASAP7_75t_R _08357_ (.A(_02519_),
    .Y(_02520_));
 INVx1_ASAP7_75t_R _08358_ (.A(_00104_),
    .Y(_02521_));
 OAI21x1_ASAP7_75t_R _08359_ (.A1(_02453_),
    .A2(_02492_),
    .B(_02521_),
    .Y(_02522_));
 AOI21x1_ASAP7_75t_R _08360_ (.A1(_00929_),
    .A2(net2718),
    .B(_00948_),
    .Y(_02523_));
 NAND2x2_ASAP7_75t_R _08361_ (.A(net5419),
    .B(_02520_),
    .Y(_02524_));
 BUFx3_ASAP7_75t_R place3027 (.A(net3026),
    .Y(net3027));
 BUFx3_ASAP7_75t_R place3012 (.A(_05148_),
    .Y(net3012));
 NAND2x1_ASAP7_75t_R _08364_ (.A(net5249),
    .B(net5050),
    .Y(_02527_));
 BUFx3_ASAP7_75t_R place3011 (.A(_06263_),
    .Y(net3011));
 BUFx3_ASAP7_75t_R place3010 (.A(_06282_),
    .Y(net3010));
 AO21x1_ASAP7_75t_R _08367_ (.A1(net2712),
    .A2(net4688),
    .B(net5249),
    .Y(_02530_));
 OAI21x1_ASAP7_75t_R _08368_ (.A1(_02527_),
    .A2(net2704),
    .B(_02530_),
    .Y(_00683_));
 INVx1_ASAP7_75t_R _08369_ (.A(_00191_),
    .Y(_02531_));
 INVx1_ASAP7_75t_R _08370_ (.A(_00194_),
    .Y(_02532_));
 INVx1_ASAP7_75t_R _08371_ (.A(_00552_),
    .Y(_02533_));
 AND3x1_ASAP7_75t_R _08372_ (.A(net4926),
    .B(net4925),
    .C(_02533_),
    .Y(_02534_));
 INVx1_ASAP7_75t_R _08373_ (.A(_00189_),
    .Y(_02535_));
 AND3x1_ASAP7_75t_R _08374_ (.A(_02534_),
    .B(net4924),
    .C(net5057),
    .Y(_02536_));
 INVx1_ASAP7_75t_R _08375_ (.A(net5225),
    .Y(_02537_));
 INVx1_ASAP7_75t_R _08376_ (.A(_00188_),
    .Y(_02538_));
 AND3x1_ASAP7_75t_R _08377_ (.A(_02536_),
    .B(_02537_),
    .C(net4922),
    .Y(_02539_));
 INVx1_ASAP7_75t_R _08378_ (.A(net5223),
    .Y(_02540_));
 INVx1_ASAP7_75t_R _08379_ (.A(net5224),
    .Y(_02541_));
 AND3x1_ASAP7_75t_R _08380_ (.A(net4576),
    .B(_02540_),
    .C(_02541_),
    .Y(_02542_));
 XNOR2x2_ASAP7_75t_R _08381_ (.A(net5248),
    .B(_02542_),
    .Y(_02543_));
 NAND2x1_ASAP7_75t_R _08382_ (.A(net5051),
    .B(_02543_),
    .Y(_02544_));
 BUFx3_ASAP7_75t_R place3009 (.A(_06294_),
    .Y(net3009));
 AO21x1_ASAP7_75t_R _08384_ (.A1(net2712),
    .A2(net4688),
    .B(net5248),
    .Y(_02546_));
 OAI21x1_ASAP7_75t_R _08385_ (.A1(_02544_),
    .A2(net2704),
    .B(_02546_),
    .Y(_00684_));
 AND3x1_ASAP7_75t_R _08386_ (.A(_02532_),
    .B(\u_hamming_window.calc_pointer[1] ),
    .C(\u_hamming_window.calc_pointer[0] ),
    .Y(_02547_));
 AND3x1_ASAP7_75t_R _08387_ (.A(_02547_),
    .B(_00922_),
    .C(_02531_),
    .Y(_02548_));
 AND3x1_ASAP7_75t_R _08388_ (.A(_02548_),
    .B(_02538_),
    .C(_02535_),
    .Y(_02549_));
 AND2x2_ASAP7_75t_R _08389_ (.A(_02549_),
    .B(_00924_),
    .Y(_02550_));
 INVx1_ASAP7_75t_R _08390_ (.A(net5248),
    .Y(_02551_));
 AND3x1_ASAP7_75t_R _08391_ (.A(net4637),
    .B(_02540_),
    .C(_02551_),
    .Y(_02552_));
 XNOR2x2_ASAP7_75t_R _08392_ (.A(net5247),
    .B(_02552_),
    .Y(_02553_));
 NAND2x1_ASAP7_75t_R _08393_ (.A(net5051),
    .B(_02553_),
    .Y(_02554_));
 AO21x1_ASAP7_75t_R _08394_ (.A1(net2712),
    .A2(net4688),
    .B(net5247),
    .Y(_02555_));
 OAI21x1_ASAP7_75t_R _08395_ (.A1(_02554_),
    .A2(net2704),
    .B(_02555_),
    .Y(_00685_));
 INVx1_ASAP7_75t_R _08396_ (.A(_02539_),
    .Y(_02556_));
 NOR2x1_ASAP7_75t_R _08397_ (.A(net5224),
    .B(_02556_),
    .Y(_02557_));
 INVx1_ASAP7_75t_R _08398_ (.A(net4471),
    .Y(_02558_));
 OR4x1_ASAP7_75t_R _08399_ (.A(_02558_),
    .B(net5223),
    .C(net5247),
    .D(net5248),
    .Y(_02559_));
 XOR2x2_ASAP7_75t_R _08400_ (.A(_02559_),
    .B(net5246),
    .Y(_02560_));
 NAND2x1_ASAP7_75t_R _08401_ (.A(net5051),
    .B(_02560_),
    .Y(_02561_));
 AO21x1_ASAP7_75t_R _08402_ (.A1(net2712),
    .A2(net4688),
    .B(net5246),
    .Y(_02562_));
 OAI21x1_ASAP7_75t_R _08403_ (.A1(_02561_),
    .A2(net5536),
    .B(_02562_),
    .Y(_00686_));
 OR4x1_ASAP7_75t_R _08404_ (.A(_00185_),
    .B(_00212_),
    .C(_00213_),
    .D(_00214_),
    .Y(_02563_));
 INVx1_ASAP7_75t_R _08405_ (.A(_02563_),
    .Y(_02564_));
 AND3x1_ASAP7_75t_R _08406_ (.A(net4686),
    .B(net5056),
    .C(net4851),
    .Y(_02565_));
 INVx1_ASAP7_75t_R _08407_ (.A(_00211_),
    .Y(_02566_));
 XOR2x2_ASAP7_75t_R _08408_ (.A(_02565_),
    .B(net4920),
    .Y(_02567_));
 NAND2x1_ASAP7_75t_R _08409_ (.A(net5052),
    .B(_02567_),
    .Y(_02568_));
 AO21x1_ASAP7_75t_R _08410_ (.A1(net4689),
    .A2(net5895),
    .B(_00211_),
    .Y(_02569_));
 OAI21x1_ASAP7_75t_R _08411_ (.A1(_02568_),
    .A2(net2705),
    .B(_02569_),
    .Y(_00687_));
 AND3x1_ASAP7_75t_R _08412_ (.A(net4471),
    .B(net4920),
    .C(net4851),
    .Y(_02570_));
 INVx1_ASAP7_75t_R _08413_ (.A(_00210_),
    .Y(_02571_));
 XOR2x2_ASAP7_75t_R _08414_ (.A(_02570_),
    .B(net4919),
    .Y(_02572_));
 NAND2x1_ASAP7_75t_R _08415_ (.A(net5052),
    .B(_02572_),
    .Y(_02573_));
 AO21x1_ASAP7_75t_R _08416_ (.A1(net4689),
    .A2(net5895),
    .B(net5245),
    .Y(_02574_));
 OAI21x1_ASAP7_75t_R _08417_ (.A1(_02573_),
    .A2(net2705),
    .B(_02574_),
    .Y(_00688_));
 AND4x1_ASAP7_75t_R _08418_ (.A(net4637),
    .B(net4919),
    .C(net4920),
    .D(net4851),
    .Y(_02575_));
 INVx1_ASAP7_75t_R _08419_ (.A(_00209_),
    .Y(_02576_));
 XOR2x2_ASAP7_75t_R _08420_ (.A(_02575_),
    .B(net4918),
    .Y(_02577_));
 NAND2x1_ASAP7_75t_R _08421_ (.A(net5052),
    .B(_02577_),
    .Y(_02578_));
 AO21x1_ASAP7_75t_R _08422_ (.A1(net2712),
    .A2(net4688),
    .B(net5244),
    .Y(_02579_));
 OAI21x1_ASAP7_75t_R _08423_ (.A1(_02578_),
    .A2(net2704),
    .B(_02579_),
    .Y(_00689_));
 AND5x1_ASAP7_75t_R _08424_ (.A(net4918),
    .B(net4471),
    .C(net4919),
    .D(net4920),
    .E(net4851),
    .Y(_02580_));
 INVx1_ASAP7_75t_R _08425_ (.A(_00208_),
    .Y(_02581_));
 XOR2x2_ASAP7_75t_R _08426_ (.A(_02580_),
    .B(_02581_),
    .Y(_02582_));
 NAND2x1_ASAP7_75t_R _08427_ (.A(net5052),
    .B(_02582_),
    .Y(_02583_));
 AO21x1_ASAP7_75t_R _08428_ (.A1(net2712),
    .A2(net4688),
    .B(net5243),
    .Y(_02584_));
 OAI21x1_ASAP7_75t_R _08429_ (.A1(_02583_),
    .A2(net5536),
    .B(_02584_),
    .Y(_00690_));
 AND5x1_ASAP7_75t_R _08430_ (.A(_02581_),
    .B(_02564_),
    .C(_02576_),
    .D(_02571_),
    .E(_02566_),
    .Y(_02585_));
 AND2x2_ASAP7_75t_R _08431_ (.A(_02585_),
    .B(_02550_),
    .Y(_02586_));
 INVx1_ASAP7_75t_R _08432_ (.A(_00207_),
    .Y(_02587_));
 XOR2x2_ASAP7_75t_R _08433_ (.A(_02586_),
    .B(net4917),
    .Y(_02588_));
 NAND2x1_ASAP7_75t_R _08434_ (.A(net5052),
    .B(_02588_),
    .Y(_02589_));
 AO21x1_ASAP7_75t_R _08435_ (.A1(net2712),
    .A2(net4688),
    .B(_00207_),
    .Y(_02590_));
 OAI21x1_ASAP7_75t_R _08436_ (.A1(_02589_),
    .A2(net2704),
    .B(_02590_),
    .Y(_00691_));
 AND3x1_ASAP7_75t_R _08437_ (.A(_02585_),
    .B(_02557_),
    .C(net4917),
    .Y(_02591_));
 INVx1_ASAP7_75t_R _08438_ (.A(_00206_),
    .Y(_02592_));
 XOR2x2_ASAP7_75t_R _08439_ (.A(net4431),
    .B(net4916),
    .Y(_02593_));
 NAND2x1_ASAP7_75t_R _08440_ (.A(net5052),
    .B(_02593_),
    .Y(_02594_));
 AO21x1_ASAP7_75t_R _08441_ (.A1(net2712),
    .A2(net4688),
    .B(_00206_),
    .Y(_02595_));
 OAI21x1_ASAP7_75t_R _08442_ (.A1(_02594_),
    .A2(net2704),
    .B(_02595_),
    .Y(_00692_));
 BUFx3_ASAP7_75t_R place3008 (.A(_06308_),
    .Y(net3008));
 BUFx3_ASAP7_75t_R place3007 (.A(_02219_),
    .Y(net3007));
 AND3x1_ASAP7_75t_R _08445_ (.A(_02586_),
    .B(_02592_),
    .C(_02587_),
    .Y(_02598_));
 INVx1_ASAP7_75t_R _08446_ (.A(net5242),
    .Y(_02599_));
 XOR2x2_ASAP7_75t_R _08447_ (.A(net4528),
    .B(net4915),
    .Y(_02600_));
 NAND2x1_ASAP7_75t_R _08448_ (.A(net5055),
    .B(_02600_),
    .Y(_02601_));
 BUFx3_ASAP7_75t_R place3005 (.A(_03925_),
    .Y(net3005));
 AO21x1_ASAP7_75t_R _08450_ (.A1(net2712),
    .A2(net4688),
    .B(net5242),
    .Y(_02603_));
 OAI21x1_ASAP7_75t_R _08451_ (.A1(_02601_),
    .A2(net5536),
    .B(_02603_),
    .Y(_00693_));
 OR2x2_ASAP7_75t_R _08452_ (.A(net5212),
    .B(_00551_),
    .Y(_02604_));
 BUFx6f_ASAP7_75t_R place3003 (.A(_03946_),
    .Y(net3003));
 AO21x1_ASAP7_75t_R _08454_ (.A1(net2712),
    .A2(net4688),
    .B(net5241),
    .Y(_02606_));
 OAI21x1_ASAP7_75t_R _08455_ (.A1(_02604_),
    .A2(net5536),
    .B(_02606_),
    .Y(_00694_));
 AND3x1_ASAP7_75t_R _08456_ (.A(_02591_),
    .B(net4915),
    .C(net4916),
    .Y(_02607_));
 INVx1_ASAP7_75t_R _08457_ (.A(_00204_),
    .Y(_02608_));
 XOR2x2_ASAP7_75t_R _08458_ (.A(_02607_),
    .B(net4914),
    .Y(_02609_));
 NAND2x1_ASAP7_75t_R _08459_ (.A(net5055),
    .B(_02609_),
    .Y(_02610_));
 AO21x1_ASAP7_75t_R _08460_ (.A1(net2713),
    .A2(net4689),
    .B(_00204_),
    .Y(_02611_));
 OAI21x1_ASAP7_75t_R _08461_ (.A1(_02610_),
    .A2(net2705),
    .B(_02611_),
    .Y(_00695_));
 AND3x1_ASAP7_75t_R _08462_ (.A(_02598_),
    .B(_02608_),
    .C(_02599_),
    .Y(_02612_));
 INVx1_ASAP7_75t_R _08463_ (.A(net5240),
    .Y(_02613_));
 XOR2x2_ASAP7_75t_R _08464_ (.A(_02612_),
    .B(net4913),
    .Y(_02614_));
 NAND2x1_ASAP7_75t_R _08465_ (.A(net5055),
    .B(_02614_),
    .Y(_02615_));
 AO21x1_ASAP7_75t_R _08466_ (.A1(net2713),
    .A2(net4689),
    .B(net5240),
    .Y(_02616_));
 OAI21x1_ASAP7_75t_R _08467_ (.A1(_02615_),
    .A2(net2705),
    .B(_02616_),
    .Y(_00696_));
 AND3x1_ASAP7_75t_R _08468_ (.A(_02607_),
    .B(net4913),
    .C(net4914),
    .Y(_02617_));
 INVx1_ASAP7_75t_R _08469_ (.A(net5239),
    .Y(_02618_));
 XOR2x2_ASAP7_75t_R _08470_ (.A(_02617_),
    .B(net4912),
    .Y(_02619_));
 NAND2x1_ASAP7_75t_R _08471_ (.A(net5055),
    .B(_02619_),
    .Y(_02620_));
 AO21x1_ASAP7_75t_R _08472_ (.A1(net2713),
    .A2(net4689),
    .B(net5239),
    .Y(_02621_));
 OAI21x1_ASAP7_75t_R _08473_ (.A1(_02620_),
    .A2(net2705),
    .B(_02621_),
    .Y(_00697_));
 AND3x1_ASAP7_75t_R _08474_ (.A(_02612_),
    .B(_02618_),
    .C(_02613_),
    .Y(_02622_));
 INVx1_ASAP7_75t_R _08475_ (.A(net5238),
    .Y(_02623_));
 XOR2x2_ASAP7_75t_R _08476_ (.A(net4430),
    .B(net4911),
    .Y(_02624_));
 NAND2x1_ASAP7_75t_R _08477_ (.A(net5055),
    .B(_02624_),
    .Y(_02625_));
 AO21x1_ASAP7_75t_R _08478_ (.A1(net2713),
    .A2(net4689),
    .B(net5238),
    .Y(_02626_));
 OAI21x1_ASAP7_75t_R _08479_ (.A1(_02625_),
    .A2(net2705),
    .B(_02626_),
    .Y(_00698_));
 AND3x1_ASAP7_75t_R _08480_ (.A(_02617_),
    .B(net4911),
    .C(net4912),
    .Y(_02627_));
 INVx1_ASAP7_75t_R _08481_ (.A(net5237),
    .Y(_02628_));
 XOR2x2_ASAP7_75t_R _08482_ (.A(_02627_),
    .B(net4910),
    .Y(_02629_));
 NAND2x1_ASAP7_75t_R _08483_ (.A(net5055),
    .B(_02629_),
    .Y(_02630_));
 AO21x1_ASAP7_75t_R _08484_ (.A1(net2713),
    .A2(net4689),
    .B(net5237),
    .Y(_02631_));
 OAI21x1_ASAP7_75t_R _08485_ (.A1(_02630_),
    .A2(net2705),
    .B(_02631_),
    .Y(_00699_));
 AND3x1_ASAP7_75t_R _08486_ (.A(_02622_),
    .B(_02628_),
    .C(_02623_),
    .Y(_02632_));
 INVx1_ASAP7_75t_R _08487_ (.A(net5236),
    .Y(_02633_));
 XOR2x2_ASAP7_75t_R _08488_ (.A(net4371),
    .B(net4909),
    .Y(_02634_));
 NAND2x1_ASAP7_75t_R _08489_ (.A(net5053),
    .B(_02634_),
    .Y(_02635_));
 AO21x1_ASAP7_75t_R _08490_ (.A1(net4689),
    .A2(net2713),
    .B(net5236),
    .Y(_02636_));
 OAI21x1_ASAP7_75t_R _08491_ (.A1(_02635_),
    .A2(net2705),
    .B(_02636_),
    .Y(_00700_));
 OR4x1_ASAP7_75t_R _08492_ (.A(net5236),
    .B(net5237),
    .C(net5238),
    .D(net5239),
    .Y(_02637_));
 INVx1_ASAP7_75t_R _08493_ (.A(_02617_),
    .Y(_02638_));
 NOR2x1_ASAP7_75t_R _08494_ (.A(_02637_),
    .B(_02638_),
    .Y(_02639_));
 INVx1_ASAP7_75t_R _08495_ (.A(net5235),
    .Y(_02640_));
 XOR2x2_ASAP7_75t_R _08496_ (.A(net4223),
    .B(net4908),
    .Y(_02641_));
 NAND2x1_ASAP7_75t_R _08497_ (.A(net5053),
    .B(_02641_),
    .Y(_02642_));
 AO21x1_ASAP7_75t_R _08498_ (.A1(net2713),
    .A2(net4689),
    .B(net5235),
    .Y(_02643_));
 OAI21x1_ASAP7_75t_R _08499_ (.A1(_02642_),
    .A2(net2705),
    .B(_02643_),
    .Y(_00701_));
 AND3x1_ASAP7_75t_R _08500_ (.A(_02632_),
    .B(_02640_),
    .C(_02633_),
    .Y(_02644_));
 INVx1_ASAP7_75t_R _08501_ (.A(net5234),
    .Y(_02645_));
 XOR2x2_ASAP7_75t_R _08502_ (.A(net4327),
    .B(net4907),
    .Y(_02646_));
 NAND2x1_ASAP7_75t_R _08503_ (.A(net5055),
    .B(_02646_),
    .Y(_02647_));
 AO21x1_ASAP7_75t_R _08504_ (.A1(net2713),
    .A2(net4689),
    .B(net5234),
    .Y(_02648_));
 OAI21x1_ASAP7_75t_R _08505_ (.A1(_02647_),
    .A2(net2705),
    .B(_02648_),
    .Y(_00702_));
 BUFx3_ASAP7_75t_R place3001 (.A(_03956_),
    .Y(net3001));
 OR4x1_ASAP7_75t_R _08507_ (.A(_02638_),
    .B(net5234),
    .C(net5235),
    .D(_02637_),
    .Y(_02650_));
 XOR2x2_ASAP7_75t_R _08508_ (.A(_02650_),
    .B(net5233),
    .Y(_02651_));
 NAND2x1_ASAP7_75t_R _08509_ (.A(net5054),
    .B(_02651_),
    .Y(_02652_));
 BUFx3_ASAP7_75t_R place3002 (.A(net3001),
    .Y(net3002));
 AO21x1_ASAP7_75t_R _08511_ (.A1(net2713),
    .A2(net4689),
    .B(net5233),
    .Y(_02654_));
 OAI21x1_ASAP7_75t_R _08512_ (.A1(_02652_),
    .A2(net2705),
    .B(_02654_),
    .Y(_00703_));
 BUFx3_ASAP7_75t_R place3004 (.A(_03943_),
    .Y(net3004));
 INVx1_ASAP7_75t_R _08514_ (.A(net5233),
    .Y(_02656_));
 AND3x1_ASAP7_75t_R _08515_ (.A(_02644_),
    .B(_02656_),
    .C(net4907),
    .Y(_02657_));
 INVx1_ASAP7_75t_R _08516_ (.A(net5232),
    .Y(_02658_));
 XOR2x2_ASAP7_75t_R _08517_ (.A(_02657_),
    .B(_02658_),
    .Y(_02659_));
 NAND2x1_ASAP7_75t_R _08518_ (.A(net5053),
    .B(_02659_),
    .Y(_02660_));
 BUFx3_ASAP7_75t_R place3000 (.A(_05159_),
    .Y(net3000));
 AO21x1_ASAP7_75t_R _08520_ (.A1(net5895),
    .A2(net4689),
    .B(net5232),
    .Y(_02662_));
 OAI21x1_ASAP7_75t_R _08521_ (.A1(_02660_),
    .A2(net2705),
    .B(_02662_),
    .Y(_00704_));
 NAND2x1_ASAP7_75t_R _08522_ (.A(net4814),
    .B(net4925),
    .Y(_02663_));
 NAND2x1_ASAP7_75t_R _08523_ (.A(net5231),
    .B(net4743),
    .Y(_02664_));
 AO21x1_ASAP7_75t_R _08524_ (.A1(_02663_),
    .A2(_02664_),
    .B(net5212),
    .Y(_02665_));
 AO21x1_ASAP7_75t_R _08525_ (.A1(net5418),
    .A2(net4688),
    .B(net5231),
    .Y(_02666_));
 OAI21x1_ASAP7_75t_R _08526_ (.A1(_02665_),
    .A2(net2704),
    .B(_02666_),
    .Y(_00705_));
 AND3x1_ASAP7_75t_R _08527_ (.A(_02658_),
    .B(_02656_),
    .C(_02645_),
    .Y(_02667_));
 AND3x1_ASAP7_75t_R _08528_ (.A(_02639_),
    .B(net4908),
    .C(_02667_),
    .Y(_02668_));
 INVx1_ASAP7_75t_R _08529_ (.A(net5230),
    .Y(_02669_));
 XOR2x2_ASAP7_75t_R _08530_ (.A(_02668_),
    .B(net4906),
    .Y(_02670_));
 NAND2x1_ASAP7_75t_R _08531_ (.A(net5053),
    .B(_02670_),
    .Y(_02671_));
 AO21x1_ASAP7_75t_R _08532_ (.A1(net5895),
    .A2(net4689),
    .B(net5230),
    .Y(_02672_));
 OAI21x1_ASAP7_75t_R _08533_ (.A1(_02671_),
    .A2(net2705),
    .B(_02672_),
    .Y(_00706_));
 AND3x1_ASAP7_75t_R _08534_ (.A(_02644_),
    .B(_02669_),
    .C(_02667_),
    .Y(_02673_));
 XNOR2x2_ASAP7_75t_R _08535_ (.A(net5229),
    .B(_02673_),
    .Y(_02674_));
 NAND2x1_ASAP7_75t_R _08536_ (.A(net5053),
    .B(_02674_),
    .Y(_02675_));
 AO21x1_ASAP7_75t_R _08537_ (.A1(net5895),
    .A2(net4689),
    .B(net5229),
    .Y(_02676_));
 OAI21x1_ASAP7_75t_R _08538_ (.A1(_02675_),
    .A2(net2705),
    .B(_02676_),
    .Y(_00707_));
 XOR2x2_ASAP7_75t_R _08539_ (.A(net4852),
    .B(net4926),
    .Y(_02677_));
 NAND2x1_ASAP7_75t_R _08540_ (.A(net5053),
    .B(_02677_),
    .Y(_02678_));
 AO21x1_ASAP7_75t_R _08541_ (.A1(net5895),
    .A2(net4689),
    .B(net5228),
    .Y(_02679_));
 OAI21x1_ASAP7_75t_R _08542_ (.A1(_02678_),
    .A2(net2705),
    .B(_02679_),
    .Y(_00708_));
 XOR2x2_ASAP7_75t_R _08543_ (.A(net4687),
    .B(net5057),
    .Y(_02680_));
 NAND2x1_ASAP7_75t_R _08544_ (.A(net5050),
    .B(_02680_),
    .Y(_02681_));
 AO21x1_ASAP7_75t_R _08545_ (.A1(net5895),
    .A2(net4689),
    .B(_00190_),
    .Y(_02682_));
 OAI21x1_ASAP7_75t_R _08546_ (.A1(_02681_),
    .A2(net2705),
    .B(_02682_),
    .Y(_00709_));
 XOR2x2_ASAP7_75t_R _08547_ (.A(net4742),
    .B(net4924),
    .Y(_02683_));
 NAND2x1_ASAP7_75t_R _08548_ (.A(net5050),
    .B(_02683_),
    .Y(_02684_));
 AO21x1_ASAP7_75t_R _08549_ (.A1(net5895),
    .A2(net4689),
    .B(net5227),
    .Y(_02685_));
 OAI21x1_ASAP7_75t_R _08550_ (.A1(_02684_),
    .A2(_02524_),
    .B(_02685_),
    .Y(_00710_));
 XOR2x2_ASAP7_75t_R _08551_ (.A(net4638),
    .B(net4922),
    .Y(_02686_));
 NAND2x1_ASAP7_75t_R _08552_ (.A(net5050),
    .B(_02686_),
    .Y(_02687_));
 AO21x1_ASAP7_75t_R _08553_ (.A1(net5895),
    .A2(net4689),
    .B(net5226),
    .Y(_02688_));
 OAI21x1_ASAP7_75t_R _08554_ (.A1(_02687_),
    .A2(net2705),
    .B(_02688_),
    .Y(_00711_));
 XOR2x2_ASAP7_75t_R _08555_ (.A(net4686),
    .B(net4923),
    .Y(_02689_));
 NAND2x1_ASAP7_75t_R _08556_ (.A(net5051),
    .B(_02689_),
    .Y(_02690_));
 AO21x1_ASAP7_75t_R _08557_ (.A1(net2712),
    .A2(net4688),
    .B(net5225),
    .Y(_02691_));
 OAI21x1_ASAP7_75t_R _08558_ (.A1(_02690_),
    .A2(net5536),
    .B(_02691_),
    .Y(_00712_));
 XOR2x2_ASAP7_75t_R _08559_ (.A(net4576),
    .B(net4921),
    .Y(_02692_));
 NAND2x1_ASAP7_75t_R _08560_ (.A(net5051),
    .B(_02692_),
    .Y(_02693_));
 AO21x1_ASAP7_75t_R _08561_ (.A1(net2712),
    .A2(net4688),
    .B(net5224),
    .Y(_02694_));
 OAI21x1_ASAP7_75t_R _08562_ (.A1(net5536),
    .A2(_02693_),
    .B(_02694_),
    .Y(_00713_));
 XOR2x2_ASAP7_75t_R _08563_ (.A(net4637),
    .B(_02540_),
    .Y(_02695_));
 NAND2x1_ASAP7_75t_R _08564_ (.A(net5051),
    .B(_02695_),
    .Y(_02696_));
 AO21x1_ASAP7_75t_R _08565_ (.A1(net2712),
    .A2(net4688),
    .B(net5223),
    .Y(_02697_));
 OAI21x1_ASAP7_75t_R _08566_ (.A1(_02696_),
    .A2(net5536),
    .B(_02697_),
    .Y(_00714_));
 BUFx3_ASAP7_75t_R place2999 (.A(_05176_),
    .Y(net2999));
 NOR2x1_ASAP7_75t_R _08568_ (.A(net5362),
    .B(net5203),
    .Y(_02699_));
 AO21x1_ASAP7_75t_R _08569_ (.A1(net5362),
    .A2(net210),
    .B(_02699_),
    .Y(_00742_));
 INVx1_ASAP7_75t_R _08570_ (.A(_00315_),
    .Y(_02700_));
 AO21x1_ASAP7_75t_R _08571_ (.A1(_02700_),
    .A2(net209),
    .B(net212),
    .Y(_02701_));
 BUFx3_ASAP7_75t_R place2998 (.A(_05181_),
    .Y(net2998));
 AO21x1_ASAP7_75t_R _08573_ (.A1(_02701_),
    .A2(_06525_),
    .B(_00958_),
    .Y(_00558_));
 INVx1_ASAP7_75t_R _08574_ (.A(_00317_),
    .Y(_02703_));
 OA21x2_ASAP7_75t_R _08575_ (.A1(_00317_),
    .A2(net5201),
    .B(net5363),
    .Y(_02704_));
 OA21x2_ASAP7_75t_R _08576_ (.A1(net5017),
    .A2(_02703_),
    .B(_02704_),
    .Y(_00557_));
 AND3x1_ASAP7_75t_R _08577_ (.A(net5041),
    .B(_02703_),
    .C(net5363),
    .Y(_00559_));
 NOR2x1p5_ASAP7_75t_R _08578_ (.A(_00161_),
    .B(_00972_),
    .Y(_02705_));
 INVx1_ASAP7_75t_R _08579_ (.A(net4636),
    .Y(_02706_));
 OA21x2_ASAP7_75t_R _08580_ (.A1(\tx_fifo.read_ptr[0] ),
    .A2(net4636),
    .B(net5362),
    .Y(_02707_));
 OA21x2_ASAP7_75t_R _08581_ (.A1(net5357),
    .A2(_02706_),
    .B(_02707_),
    .Y(_00560_));
 AO21x1_ASAP7_75t_R _08582_ (.A1(_00546_),
    .A2(net4636),
    .B(net5361),
    .Y(_02708_));
 AOI21x1_ASAP7_75t_R _08583_ (.A1(net5356),
    .A2(net4575),
    .B(_02708_),
    .Y(_00561_));
 INVx1_ASAP7_75t_R _08584_ (.A(net5355),
    .Y(_02709_));
 INVx1_ASAP7_75t_R _08585_ (.A(_00547_),
    .Y(_02710_));
 AND3x1_ASAP7_75t_R _08586_ (.A(_02710_),
    .B(net4905),
    .C(_02705_),
    .Y(_02711_));
 INVx1_ASAP7_75t_R _08587_ (.A(net4574),
    .Y(_02712_));
 AO21x1_ASAP7_75t_R _08588_ (.A1(net4636),
    .A2(_02710_),
    .B(net4905),
    .Y(_02713_));
 AND3x1_ASAP7_75t_R _08589_ (.A(_02712_),
    .B(net5362),
    .C(_02713_),
    .Y(_00562_));
 INVx1_ASAP7_75t_R _08590_ (.A(net5354),
    .Y(_02714_));
 AND3x1_ASAP7_75t_R _08591_ (.A(net4905),
    .B(\tx_fifo.read_ptr[1] ),
    .C(\tx_fifo.read_ptr[0] ),
    .Y(_02715_));
 AND3x1_ASAP7_75t_R _08592_ (.A(_02715_),
    .B(_02714_),
    .C(_02705_),
    .Y(_02716_));
 INVx1_ASAP7_75t_R _08593_ (.A(_02716_),
    .Y(_02717_));
 AO21x1_ASAP7_75t_R _08594_ (.A1(_02705_),
    .A2(_02715_),
    .B(net4904),
    .Y(_02718_));
 AND3x1_ASAP7_75t_R _08595_ (.A(_02717_),
    .B(net5362),
    .C(_02718_),
    .Y(_00563_));
 INVx1_ASAP7_75t_R _08596_ (.A(net5353),
    .Y(_02719_));
 AND3x1_ASAP7_75t_R _08597_ (.A(_02711_),
    .B(_02719_),
    .C(net4904),
    .Y(_02720_));
 INVx1_ASAP7_75t_R _08598_ (.A(_02720_),
    .Y(_02721_));
 AO21x1_ASAP7_75t_R _08599_ (.A1(net4574),
    .A2(net4904),
    .B(_02719_),
    .Y(_02722_));
 AND3x1_ASAP7_75t_R _08600_ (.A(_02721_),
    .B(net5362),
    .C(_02722_),
    .Y(_00564_));
 INVx1_ASAP7_75t_R _08601_ (.A(net5352),
    .Y(_02723_));
 AND3x1_ASAP7_75t_R _08602_ (.A(_02723_),
    .B(_02716_),
    .C(_02719_),
    .Y(_02724_));
 INVx2_ASAP7_75t_R _08603_ (.A(_02724_),
    .Y(_02725_));
 AO21x1_ASAP7_75t_R _08604_ (.A1(_02716_),
    .A2(_02719_),
    .B(_02723_),
    .Y(_02726_));
 AND3x1_ASAP7_75t_R _08605_ (.A(_02725_),
    .B(net5362),
    .C(_02726_),
    .Y(_00565_));
 OR3x1_ASAP7_75t_R _08606_ (.A(_02721_),
    .B(net5351),
    .C(net5352),
    .Y(_02727_));
 OAI21x1_ASAP7_75t_R _08607_ (.A1(net5352),
    .A2(_02721_),
    .B(net5351),
    .Y(_02728_));
 AND3x1_ASAP7_75t_R _08608_ (.A(_02727_),
    .B(net5362),
    .C(_02728_),
    .Y(_00566_));
 OR3x1_ASAP7_75t_R _08609_ (.A(_02725_),
    .B(net5350),
    .C(net5351),
    .Y(_02729_));
 OAI21x1_ASAP7_75t_R _08610_ (.A1(_02725_),
    .A2(net5351),
    .B(net5350),
    .Y(_02730_));
 AND3x1_ASAP7_75t_R _08611_ (.A(_02730_),
    .B(net5362),
    .C(_02729_),
    .Y(_00567_));
 INVx1_ASAP7_75t_R _08612_ (.A(_00307_),
    .Y(_02731_));
 AND3x1_ASAP7_75t_R _08613_ (.A(_02731_),
    .B(net5039),
    .C(net5040),
    .Y(_02732_));
 INVx1_ASAP7_75t_R _08614_ (.A(_00305_),
    .Y(_02733_));
 INVx1_ASAP7_75t_R _08615_ (.A(net5346),
    .Y(_02734_));
 AND3x1_ASAP7_75t_R _08616_ (.A(_02732_),
    .B(_02733_),
    .C(_02734_),
    .Y(_02735_));
 XNOR2x2_ASAP7_75t_R _08617_ (.A(net5036),
    .B(net4741),
    .Y(_02736_));
 INVx1_ASAP7_75t_R _08618_ (.A(net5344),
    .Y(_02737_));
 OR3x1_ASAP7_75t_R _08619_ (.A(_00468_),
    .B(_00307_),
    .C(_00306_),
    .Y(_02738_));
 INVx1_ASAP7_75t_R _08620_ (.A(_02738_),
    .Y(_02739_));
 NAND2x1_ASAP7_75t_R _08621_ (.A(_02739_),
    .B(_02733_),
    .Y(_02740_));
 NOR2x1_ASAP7_75t_R _08622_ (.A(net5345),
    .B(_02740_),
    .Y(_02741_));
 NAND2x1_ASAP7_75t_R _08623_ (.A(_02741_),
    .B(_02737_),
    .Y(_02742_));
 NOR2x1_ASAP7_75t_R _08624_ (.A(net5343),
    .B(_02742_),
    .Y(_02743_));
 XOR2x2_ASAP7_75t_R _08625_ (.A(_00307_),
    .B(net4822),
    .Y(_02744_));
 XOR2x2_ASAP7_75t_R _08626_ (.A(_02744_),
    .B(_02709_),
    .Y(_02745_));
 XOR2x2_ASAP7_75t_R _08627_ (.A(net4759),
    .B(net5356),
    .Y(_02746_));
 OR4x1_ASAP7_75t_R _08628_ (.A(_02743_),
    .B(_00970_),
    .C(_02745_),
    .D(_02746_),
    .Y(_02747_));
 XOR2x2_ASAP7_75t_R _08629_ (.A(net4573),
    .B(net5037),
    .Y(_02748_));
 XOR2x2_ASAP7_75t_R _08630_ (.A(net4850),
    .B(net4903),
    .Y(_02749_));
 XNOR2x2_ASAP7_75t_R _08631_ (.A(_00965_),
    .B(net4740),
    .Y(_02750_));
 OAI21x1_ASAP7_75t_R _08632_ (.A1(net5354),
    .A2(_02749_),
    .B(_02750_),
    .Y(_02751_));
 AO21x1_ASAP7_75t_R _08633_ (.A1(net5354),
    .A2(_02749_),
    .B(_02751_),
    .Y(_02752_));
 INVx1_ASAP7_75t_R _08634_ (.A(net5345),
    .Y(_02753_));
 AND3x1_ASAP7_75t_R _08635_ (.A(_02735_),
    .B(_02737_),
    .C(_02753_),
    .Y(_02754_));
 XOR2x2_ASAP7_75t_R _08636_ (.A(_02754_),
    .B(net5038),
    .Y(_02755_));
 OR5x1_ASAP7_75t_R _08637_ (.A(_02747_),
    .B(_02736_),
    .C(_02748_),
    .D(_02752_),
    .E(_02755_),
    .Y(_02756_));
 INVx1_ASAP7_75t_R _08638_ (.A(_00545_),
    .Y(_02757_));
 AND4x1_ASAP7_75t_R _08639_ (.A(net5350),
    .B(net5351),
    .C(net5352),
    .D(net5353),
    .Y(_02758_));
 AND5x1_ASAP7_75t_R _08640_ (.A(net5354),
    .B(_02743_),
    .C(net5355),
    .D(_02757_),
    .E(_02758_),
    .Y(_02759_));
 NOR2x1_ASAP7_75t_R _08641_ (.A(_00333_),
    .B(_02759_),
    .Y(_02760_));
 AND2x4_ASAP7_75t_R _08642_ (.A(_02760_),
    .B(_02756_),
    .Y(_02761_));
 INVx4_ASAP7_75t_R _08643_ (.A(net4326),
    .Y(_02762_));
 OA21x2_ASAP7_75t_R _08644_ (.A1(net4326),
    .A2(net5040),
    .B(net5362),
    .Y(_02763_));
 OA21x2_ASAP7_75t_R _08645_ (.A1(net5349),
    .A2(_02762_),
    .B(_02763_),
    .Y(_00568_));
 AO21x1_ASAP7_75t_R _08646_ (.A1(net4326),
    .A2(net4759),
    .B(net5361),
    .Y(_02764_));
 AOI21x1_ASAP7_75t_R _08647_ (.A1(net5348),
    .A2(net4279),
    .B(_02764_),
    .Y(_00569_));
 OA21x2_ASAP7_75t_R _08648_ (.A1(net4326),
    .A2(_02731_),
    .B(net5362),
    .Y(_02765_));
 OA21x2_ASAP7_75t_R _08649_ (.A1(_02744_),
    .A2(_02762_),
    .B(_02765_),
    .Y(_00570_));
 OA21x2_ASAP7_75t_R _08650_ (.A1(net4326),
    .A2(net4903),
    .B(net5362),
    .Y(_02766_));
 OA21x2_ASAP7_75t_R _08651_ (.A1(_02749_),
    .A2(_02762_),
    .B(_02766_),
    .Y(_00571_));
 AO21x1_ASAP7_75t_R _08652_ (.A1(_02739_),
    .A2(net4326),
    .B(_02733_),
    .Y(_02767_));
 OA211x2_ASAP7_75t_R _08653_ (.A1(_02740_),
    .A2(_02762_),
    .B(_02767_),
    .C(net5362),
    .Y(_00572_));
 AND3x1_ASAP7_75t_R _08654_ (.A(_02761_),
    .B(net4902),
    .C(net4741),
    .Y(_02768_));
 INVx1_ASAP7_75t_R _08655_ (.A(_02768_),
    .Y(_02769_));
 AO21x1_ASAP7_75t_R _08656_ (.A1(net4326),
    .A2(net4741),
    .B(net4902),
    .Y(_02770_));
 AND3x1_ASAP7_75t_R _08657_ (.A(_02769_),
    .B(net5362),
    .C(_02770_),
    .Y(_00573_));
 AO21x1_ASAP7_75t_R _08658_ (.A1(net4573),
    .A2(net4326),
    .B(_02737_),
    .Y(_02771_));
 OA211x2_ASAP7_75t_R _08659_ (.A1(_02742_),
    .A2(_02762_),
    .B(_02771_),
    .C(net5362),
    .Y(_00574_));
 OR3x1_ASAP7_75t_R _08660_ (.A(_02769_),
    .B(net5343),
    .C(net5344),
    .Y(_02772_));
 OAI21x1_ASAP7_75t_R _08661_ (.A1(net5344),
    .A2(net4222),
    .B(net5343),
    .Y(_02773_));
 AND3x1_ASAP7_75t_R _08662_ (.A(_02772_),
    .B(net5362),
    .C(_02773_),
    .Y(_00575_));
 NOR2x1_ASAP7_75t_R _08663_ (.A(net5340),
    .B(net5361),
    .Y(_00576_));
 NOR2x1_ASAP7_75t_R _08664_ (.A(net5342),
    .B(net4861),
    .Y(_02774_));
 AO21x2_ASAP7_75t_R _08665_ (.A1(_00319_),
    .A2(_00942_),
    .B(_00938_),
    .Y(_02775_));
 INVx3_ASAP7_75t_R _08666_ (.A(net4849),
    .Y(_02776_));
 OA21x2_ASAP7_75t_R _08667_ (.A1(_02776_),
    .A2(_00470_),
    .B(net5362),
    .Y(_02777_));
 OA21x2_ASAP7_75t_R _08668_ (.A1(\u_dct.k_ptr[0] ),
    .A2(_02774_),
    .B(_02777_),
    .Y(_00577_));
 NOR2x1_ASAP7_75t_R _08669_ (.A(_00473_),
    .B(net5361),
    .Y(_02778_));
 AO32x1_ASAP7_75t_R _08670_ (.A1(net5362),
    .A2(\u_dct.k_ptr[1] ),
    .A3(_02776_),
    .B1(_02774_),
    .B2(_02778_),
    .Y(_00578_));
 OR3x1_ASAP7_75t_R _08671_ (.A(_02776_),
    .B(_00474_),
    .C(net5339),
    .Y(_02779_));
 OAI21x1_ASAP7_75t_R _08672_ (.A1(_00474_),
    .A2(_02776_),
    .B(net5339),
    .Y(_02780_));
 AOI21x1_ASAP7_75t_R _08673_ (.A1(net5342),
    .A2(net5046),
    .B(net5361),
    .Y(_02781_));
 AND3x1_ASAP7_75t_R _08674_ (.A(_02779_),
    .B(_02780_),
    .C(_02781_),
    .Y(_00579_));
 OR3x1_ASAP7_75t_R _08675_ (.A(_00300_),
    .B(_00471_),
    .C(_00470_),
    .Y(_02782_));
 OR3x1_ASAP7_75t_R _08676_ (.A(_02776_),
    .B(net5338),
    .C(_02782_),
    .Y(_02783_));
 OAI21x1_ASAP7_75t_R _08677_ (.A1(_02782_),
    .A2(net4739),
    .B(net5338),
    .Y(_02784_));
 AND3x1_ASAP7_75t_R _08678_ (.A(_02783_),
    .B(_02781_),
    .C(_02784_),
    .Y(_00580_));
 NOR2x1p5_ASAP7_75t_R _08679_ (.A(_00321_),
    .B(_00945_),
    .Y(_02785_));
 NOR2x1p5_ASAP7_75t_R _08680_ (.A(_02785_),
    .B(_02775_),
    .Y(_02786_));
 OA21x2_ASAP7_75t_R _08681_ (.A1(net4738),
    .A2(net5002),
    .B(net5362),
    .Y(_02787_));
 OA21x2_ASAP7_75t_R _08682_ (.A1(net5337),
    .A2(net4685),
    .B(_02787_),
    .Y(_00581_));
 OR3x1_ASAP7_75t_R _08683_ (.A(net4861),
    .B(_00478_),
    .C(net5341),
    .Y(_02788_));
 NAND2x1p5_ASAP7_75t_R _08684_ (.A(net4685),
    .B(net5001),
    .Y(_02789_));
 AOI21x1_ASAP7_75t_R _08685_ (.A1(_02789_),
    .A2(_02788_),
    .B(net5361),
    .Y(_00582_));
 INVx2_ASAP7_75t_R _08686_ (.A(net4685),
    .Y(_02790_));
 INVx1_ASAP7_75t_R _08687_ (.A(_00479_),
    .Y(_02791_));
 AND3x1_ASAP7_75t_R _08688_ (.A(_02790_),
    .B(_00935_),
    .C(_02791_),
    .Y(_02792_));
 INVx2_ASAP7_75t_R _08689_ (.A(_02792_),
    .Y(_02793_));
 OA21x2_ASAP7_75t_R _08690_ (.A1(_02776_),
    .A2(_00937_),
    .B(net5362),
    .Y(_02794_));
 AO21x1_ASAP7_75t_R _08691_ (.A1(_02790_),
    .A2(_02791_),
    .B(_00935_),
    .Y(_02795_));
 AND3x1_ASAP7_75t_R _08692_ (.A(_02793_),
    .B(_02794_),
    .C(_02795_),
    .Y(_00583_));
 OR4x1_ASAP7_75t_R _08693_ (.A(_02786_),
    .B(_00298_),
    .C(_00476_),
    .D(_00475_),
    .Y(_02796_));
 NOR2x1_ASAP7_75t_R _08694_ (.A(net5335),
    .B(_02796_),
    .Y(_02797_));
 INVx1_ASAP7_75t_R _08695_ (.A(_02797_),
    .Y(_02798_));
 NAND2x1_ASAP7_75t_R _08696_ (.A(net5335),
    .B(_02796_),
    .Y(_02799_));
 AND3x1_ASAP7_75t_R _08697_ (.A(_02798_),
    .B(_02794_),
    .C(_02799_),
    .Y(_00584_));
 OR3x1_ASAP7_75t_R _08698_ (.A(_02793_),
    .B(net5334),
    .C(net5335),
    .Y(_02800_));
 OAI21x1_ASAP7_75t_R _08699_ (.A1(_02793_),
    .A2(net5335),
    .B(net5334),
    .Y(_02801_));
 AND3x1_ASAP7_75t_R _08700_ (.A(_02801_),
    .B(_02794_),
    .C(_02800_),
    .Y(_00585_));
 OR3x1_ASAP7_75t_R _08701_ (.A(_02798_),
    .B(net5333),
    .C(net5334),
    .Y(_02802_));
 OAI21x1_ASAP7_75t_R _08702_ (.A1(net5334),
    .A2(_02798_),
    .B(net5333),
    .Y(_02803_));
 AND3x1_ASAP7_75t_R _08703_ (.A(_02802_),
    .B(_02794_),
    .C(_02803_),
    .Y(_00586_));
 NOR2x1_ASAP7_75t_R _08704_ (.A(net5328),
    .B(net5361),
    .Y(_00587_));
 AO21x2_ASAP7_75t_R _08705_ (.A1(_01099_),
    .A2(_01118_),
    .B(net5329),
    .Y(_02804_));
 AOI211x1_ASAP7_75t_R _08706_ (.A1(_01131_),
    .A2(_02518_),
    .B(_01124_),
    .C(_01105_),
    .Y(_02805_));
 AND2x4_ASAP7_75t_R _08707_ (.A(_02804_),
    .B(_02805_),
    .Y(_02806_));
 AO21x2_ASAP7_75t_R _08708_ (.A1(net5331),
    .A2(net4087),
    .B(net5361),
    .Y(_02807_));
 XOR2x2_ASAP7_75t_R _08709_ (.A(net4087),
    .B(net5327),
    .Y(_02808_));
 NOR2x1_ASAP7_75t_R _08710_ (.A(_02808_),
    .B(net4045),
    .Y(_00588_));
 INVx3_ASAP7_75t_R _08711_ (.A(_02807_),
    .Y(_02809_));
 NAND2x1_ASAP7_75t_R _08712_ (.A(_00515_),
    .B(net4087),
    .Y(_02810_));
 OA211x2_ASAP7_75t_R _08713_ (.A1(\u_fft.power_ptr[1] ),
    .A2(net4087),
    .B(_02810_),
    .C(_02809_),
    .Y(_00589_));
 INVx3_ASAP7_75t_R _08714_ (.A(_02806_),
    .Y(_02811_));
 OR3x1_ASAP7_75t_R _08715_ (.A(_02811_),
    .B(net5325),
    .C(_00514_),
    .Y(_02812_));
 OAI21x1_ASAP7_75t_R _08716_ (.A1(net4821),
    .A2(net4044),
    .B(net5325),
    .Y(_02813_));
 AND3x1_ASAP7_75t_R _08717_ (.A(net4019),
    .B(net4020),
    .C(_02813_),
    .Y(_00590_));
 INVx1_ASAP7_75t_R _08718_ (.A(_00291_),
    .Y(_02814_));
 AND3x1_ASAP7_75t_R _08719_ (.A(_02814_),
    .B(\u_fft.power_ptr[1] ),
    .C(\u_fft.power_ptr[0] ),
    .Y(_02815_));
 AND3x1_ASAP7_75t_R _08720_ (.A(net4151),
    .B(net4684),
    .C(net4848),
    .Y(_02816_));
 XOR2x2_ASAP7_75t_R _08721_ (.A(_02816_),
    .B(net5324),
    .Y(_02817_));
 NOR2x1_ASAP7_75t_R _08722_ (.A(_02817_),
    .B(net4045),
    .Y(_00591_));
 NOR2x1_ASAP7_75t_R _08723_ (.A(_02812_),
    .B(net5324),
    .Y(_02818_));
 XOR2x2_ASAP7_75t_R _08724_ (.A(net4000),
    .B(net5323),
    .Y(_02819_));
 NOR2x1_ASAP7_75t_R _08725_ (.A(net4045),
    .B(_02819_),
    .Y(_00592_));
 INVx1_ASAP7_75t_R _08726_ (.A(_00289_),
    .Y(_02820_));
 INVx1_ASAP7_75t_R _08727_ (.A(_00290_),
    .Y(_02821_));
 AND3x1_ASAP7_75t_R _08728_ (.A(net4848),
    .B(_02820_),
    .C(_02821_),
    .Y(_02822_));
 INVx1_ASAP7_75t_R _08729_ (.A(_02822_),
    .Y(_02823_));
 OR3x1_ASAP7_75t_R _08730_ (.A(net4044),
    .B(net5322),
    .C(_02823_),
    .Y(_02824_));
 INVx1_ASAP7_75t_R _08731_ (.A(_00288_),
    .Y(_02825_));
 AO21x1_ASAP7_75t_R _08732_ (.A1(net4087),
    .A2(_02822_),
    .B(_02825_),
    .Y(_02826_));
 AND3x1_ASAP7_75t_R _08733_ (.A(net4020),
    .B(_02824_),
    .C(_02826_),
    .Y(_00593_));
 INVx1_ASAP7_75t_R _08734_ (.A(_00287_),
    .Y(_02827_));
 AND3x1_ASAP7_75t_R _08735_ (.A(_02820_),
    .B(_02825_),
    .C(_02818_),
    .Y(_02828_));
 INVx2_ASAP7_75t_R _08736_ (.A(_02828_),
    .Y(_02829_));
 OA21x2_ASAP7_75t_R _08737_ (.A1(_02829_),
    .A2(net5321),
    .B(_02809_),
    .Y(_02830_));
 OA21x2_ASAP7_75t_R _08738_ (.A1(net4901),
    .A2(_02828_),
    .B(_02830_),
    .Y(_00594_));
 INVx1_ASAP7_75t_R _08739_ (.A(_00286_),
    .Y(_02831_));
 AND5x1_ASAP7_75t_R _08740_ (.A(_02827_),
    .B(_02815_),
    .C(_02825_),
    .D(_02820_),
    .E(_02821_),
    .Y(_02832_));
 AND3x1_ASAP7_75t_R _08741_ (.A(net4087),
    .B(_02831_),
    .C(_02832_),
    .Y(_02833_));
 INVx2_ASAP7_75t_R _08742_ (.A(_02833_),
    .Y(_02834_));
 AO21x1_ASAP7_75t_R _08743_ (.A1(net4087),
    .A2(_02832_),
    .B(_02831_),
    .Y(_02835_));
 AND3x1_ASAP7_75t_R _08744_ (.A(_02834_),
    .B(_02835_),
    .C(net4021),
    .Y(_00595_));
 NAND2x1_ASAP7_75t_R _08745_ (.A(_02831_),
    .B(net4901),
    .Y(_02836_));
 OR3x1_ASAP7_75t_R _08746_ (.A(_02829_),
    .B(_00285_),
    .C(_02836_),
    .Y(_02837_));
 OAI21x1_ASAP7_75t_R _08747_ (.A1(_02829_),
    .A2(_02836_),
    .B(_00285_),
    .Y(_02838_));
 AND3x1_ASAP7_75t_R _08748_ (.A(_02837_),
    .B(net4021),
    .C(_02838_),
    .Y(_00596_));
 OR3x1_ASAP7_75t_R _08749_ (.A(_02834_),
    .B(_00284_),
    .C(_00285_),
    .Y(_02839_));
 OAI21x1_ASAP7_75t_R _08750_ (.A1(_02834_),
    .A2(_00285_),
    .B(_00284_),
    .Y(_02840_));
 AND3x1_ASAP7_75t_R _08751_ (.A(_02839_),
    .B(_02840_),
    .C(net4021),
    .Y(_00597_));
 INVx2_ASAP7_75t_R _08752_ (.A(_01132_),
    .Y(_02841_));
 BUFx3_ASAP7_75t_R place2997 (.A(_06309_),
    .Y(net2997));
 AO21x1_ASAP7_75t_R _08754_ (.A1(net4696),
    .A2(net5327),
    .B(net5361),
    .Y(_02843_));
 AOI21x1_ASAP7_75t_R _08755_ (.A1(net5319),
    .A2(net4634),
    .B(_02843_),
    .Y(_00598_));
 AO21x1_ASAP7_75t_R _08756_ (.A1(net5326),
    .A2(net4692),
    .B(net5361),
    .Y(_02844_));
 AOI21x1_ASAP7_75t_R _08757_ (.A1(net5318),
    .A2(net4634),
    .B(_02844_),
    .Y(_00599_));
 AO21x1_ASAP7_75t_R _08758_ (.A1(net4692),
    .A2(net5325),
    .B(net5361),
    .Y(_02845_));
 AOI21x1_ASAP7_75t_R _08759_ (.A1(net5317),
    .A2(net4633),
    .B(_02845_),
    .Y(_00600_));
 AO21x1_ASAP7_75t_R _08760_ (.A1(net4696),
    .A2(net5324),
    .B(net5361),
    .Y(_02846_));
 AOI21x1_ASAP7_75t_R _08761_ (.A1(net5316),
    .A2(net4634),
    .B(_02846_),
    .Y(_00601_));
 AO21x1_ASAP7_75t_R _08762_ (.A1(net4692),
    .A2(net5323),
    .B(net5361),
    .Y(_02847_));
 AOI21x1_ASAP7_75t_R _08763_ (.A1(net5315),
    .A2(net4633),
    .B(_02847_),
    .Y(_00602_));
 BUFx3_ASAP7_75t_R place2996 (.A(_02220_),
    .Y(net2996));
 AO21x1_ASAP7_75t_R _08765_ (.A1(net4692),
    .A2(net5322),
    .B(net5361),
    .Y(_02849_));
 AOI21x1_ASAP7_75t_R _08766_ (.A1(net5314),
    .A2(net4630),
    .B(_02849_),
    .Y(_00603_));
 AO21x1_ASAP7_75t_R _08767_ (.A1(net4692),
    .A2(net5321),
    .B(net5361),
    .Y(_02850_));
 AOI21x1_ASAP7_75t_R _08768_ (.A1(net5313),
    .A2(net4630),
    .B(_02850_),
    .Y(_00604_));
 AO21x1_ASAP7_75t_R _08769_ (.A1(net5320),
    .A2(net4692),
    .B(net5361),
    .Y(_02851_));
 AOI21x1_ASAP7_75t_R _08770_ (.A1(net5312),
    .A2(net4630),
    .B(_02851_),
    .Y(_00605_));
 BUFx3_ASAP7_75t_R place2995 (.A(_03947_),
    .Y(net2995));
 AO21x1_ASAP7_75t_R _08772_ (.A1(net4692),
    .A2(_00285_),
    .B(net5361),
    .Y(_02853_));
 AOI21x1_ASAP7_75t_R _08773_ (.A1(net5311),
    .A2(net4630),
    .B(_02853_),
    .Y(_00606_));
 AO21x1_ASAP7_75t_R _08774_ (.A1(net4692),
    .A2(_00284_),
    .B(net5361),
    .Y(_02854_));
 AOI21x1_ASAP7_75t_R _08775_ (.A1(net5310),
    .A2(net4630),
    .B(_02854_),
    .Y(_00607_));
 BUFx3_ASAP7_75t_R place2994 (.A(_03974_),
    .Y(net2994));
 AO21x1_ASAP7_75t_R _08777_ (.A1(net4696),
    .A2(_00283_),
    .B(net5361),
    .Y(_02856_));
 AOI21x1_ASAP7_75t_R _08778_ (.A1(net5309),
    .A2(net4634),
    .B(_02856_),
    .Y(_00608_));
 AO21x1_ASAP7_75t_R _08779_ (.A1(net4695),
    .A2(_00282_),
    .B(net5361),
    .Y(_02857_));
 AOI21x1_ASAP7_75t_R _08780_ (.A1(net5308),
    .A2(net4635),
    .B(_02857_),
    .Y(_00609_));
 AO21x1_ASAP7_75t_R _08781_ (.A1(net4695),
    .A2(_00281_),
    .B(net5361),
    .Y(_02858_));
 AOI21x1_ASAP7_75t_R _08782_ (.A1(net5307),
    .A2(net4635),
    .B(_02858_),
    .Y(_00610_));
 AO21x1_ASAP7_75t_R _08783_ (.A1(net4696),
    .A2(_00280_),
    .B(net5361),
    .Y(_02859_));
 AOI21x1_ASAP7_75t_R _08784_ (.A1(net5306),
    .A2(net4634),
    .B(_02859_),
    .Y(_00611_));
 AO21x1_ASAP7_75t_R _08785_ (.A1(net4695),
    .A2(_00279_),
    .B(net5361),
    .Y(_02860_));
 AOI21x1_ASAP7_75t_R _08786_ (.A1(net5305),
    .A2(net4632),
    .B(_02860_),
    .Y(_00612_));
 BUFx3_ASAP7_75t_R place2993 (.A(_05150_),
    .Y(net2993));
 AO21x1_ASAP7_75t_R _08788_ (.A1(net4693),
    .A2(_00278_),
    .B(net5361),
    .Y(_02862_));
 AOI21x1_ASAP7_75t_R _08789_ (.A1(net5304),
    .A2(net4631),
    .B(_02862_),
    .Y(_00613_));
 AO21x1_ASAP7_75t_R _08790_ (.A1(net4693),
    .A2(_00277_),
    .B(net5361),
    .Y(_02863_));
 AOI21x1_ASAP7_75t_R _08791_ (.A1(net5303),
    .A2(net4630),
    .B(_02863_),
    .Y(_00614_));
 AO21x1_ASAP7_75t_R _08792_ (.A1(net4693),
    .A2(_00276_),
    .B(net5361),
    .Y(_02864_));
 AOI21x1_ASAP7_75t_R _08793_ (.A1(net5302),
    .A2(net4630),
    .B(_02864_),
    .Y(_00615_));
 BUFx3_ASAP7_75t_R place2992 (.A(_05160_),
    .Y(net2992));
 AO21x1_ASAP7_75t_R _08795_ (.A1(net4693),
    .A2(_00275_),
    .B(net5361),
    .Y(_02866_));
 AOI21x1_ASAP7_75t_R _08796_ (.A1(net5301),
    .A2(net4630),
    .B(_02866_),
    .Y(_00616_));
 AO21x1_ASAP7_75t_R _08797_ (.A1(net4693),
    .A2(_00274_),
    .B(net5361),
    .Y(_02867_));
 AOI21x1_ASAP7_75t_R _08798_ (.A1(net5300),
    .A2(net4630),
    .B(_02867_),
    .Y(_00617_));
 BUFx3_ASAP7_75t_R place2991 (.A(_05169_),
    .Y(net2991));
 AO21x1_ASAP7_75t_R _08800_ (.A1(net4696),
    .A2(_00273_),
    .B(net5361),
    .Y(_02869_));
 AOI21x1_ASAP7_75t_R _08801_ (.A1(net5299),
    .A2(net4634),
    .B(_02869_),
    .Y(_00618_));
 AO21x1_ASAP7_75t_R _08802_ (.A1(net4695),
    .A2(_00272_),
    .B(net5361),
    .Y(_02870_));
 AOI21x1_ASAP7_75t_R _08803_ (.A1(net5298),
    .A2(net4635),
    .B(_02870_),
    .Y(_00619_));
 AO21x1_ASAP7_75t_R _08804_ (.A1(net4695),
    .A2(_00271_),
    .B(net5361),
    .Y(_02871_));
 AOI21x1_ASAP7_75t_R _08805_ (.A1(_00261_),
    .A2(net4635),
    .B(_02871_),
    .Y(_00620_));
 AO21x1_ASAP7_75t_R _08806_ (.A1(net4696),
    .A2(_00270_),
    .B(net5361),
    .Y(_02872_));
 AOI21x1_ASAP7_75t_R _08807_ (.A1(net5297),
    .A2(net4634),
    .B(_02872_),
    .Y(_00621_));
 AO21x1_ASAP7_75t_R _08808_ (.A1(net4695),
    .A2(_00269_),
    .B(net5361),
    .Y(_02873_));
 AOI21x1_ASAP7_75t_R _08809_ (.A1(net5296),
    .A2(net4632),
    .B(_02873_),
    .Y(_00622_));
 BUFx3_ASAP7_75t_R place2990 (.A(_05177_),
    .Y(net2990));
 AO21x1_ASAP7_75t_R _08811_ (.A1(net4693),
    .A2(_00268_),
    .B(net5361),
    .Y(_02875_));
 AOI21x1_ASAP7_75t_R _08812_ (.A1(_00258_),
    .A2(net4631),
    .B(_02875_),
    .Y(_00623_));
 AO21x1_ASAP7_75t_R _08813_ (.A1(net4693),
    .A2(_00267_),
    .B(net5361),
    .Y(_02876_));
 AOI21x1_ASAP7_75t_R _08814_ (.A1(net5295),
    .A2(net4630),
    .B(_02876_),
    .Y(_00624_));
 AO21x1_ASAP7_75t_R _08815_ (.A1(net4693),
    .A2(_00266_),
    .B(net5361),
    .Y(_02877_));
 AOI21x1_ASAP7_75t_R _08816_ (.A1(net5294),
    .A2(net4630),
    .B(_02877_),
    .Y(_00625_));
 BUFx3_ASAP7_75t_R place3006 (.A(net3005),
    .Y(net3006));
 AO21x1_ASAP7_75t_R _08818_ (.A1(net4693),
    .A2(_00265_),
    .B(net5361),
    .Y(_02879_));
 AOI21x1_ASAP7_75t_R _08819_ (.A1(net5293),
    .A2(net4631),
    .B(_02879_),
    .Y(_00626_));
 AO21x1_ASAP7_75t_R _08820_ (.A1(net4695),
    .A2(_00264_),
    .B(net5361),
    .Y(_02880_));
 AOI21x1_ASAP7_75t_R _08821_ (.A1(net5292),
    .A2(net4632),
    .B(_02880_),
    .Y(_00627_));
 BUFx3_ASAP7_75t_R place2988 (.A(_05182_),
    .Y(net2988));
 AO21x1_ASAP7_75t_R _08823_ (.A1(net4696),
    .A2(_00263_),
    .B(net5361),
    .Y(_02882_));
 AOI21x1_ASAP7_75t_R _08824_ (.A1(net5291),
    .A2(net4635),
    .B(_02882_),
    .Y(_00628_));
 AO21x1_ASAP7_75t_R _08825_ (.A1(net4695),
    .A2(_00262_),
    .B(net5361),
    .Y(_02883_));
 AOI21x1_ASAP7_75t_R _08826_ (.A1(net5290),
    .A2(net4635),
    .B(_02883_),
    .Y(_00629_));
 AO21x1_ASAP7_75t_R _08827_ (.A1(net4695),
    .A2(_00261_),
    .B(net5361),
    .Y(_02884_));
 AOI21x1_ASAP7_75t_R _08828_ (.A1(net5289),
    .A2(net4635),
    .B(_02884_),
    .Y(_00630_));
 AO21x1_ASAP7_75t_R _08829_ (.A1(net4696),
    .A2(_00260_),
    .B(net5361),
    .Y(_02885_));
 AOI21x1_ASAP7_75t_R _08830_ (.A1(net5288),
    .A2(net4635),
    .B(_02885_),
    .Y(_00631_));
 AO21x1_ASAP7_75t_R _08831_ (.A1(net4695),
    .A2(_00259_),
    .B(net5361),
    .Y(_02886_));
 AOI21x1_ASAP7_75t_R _08832_ (.A1(net5287),
    .A2(net4632),
    .B(_02886_),
    .Y(_00632_));
 BUFx3_ASAP7_75t_R place2987 (.A(_05191_),
    .Y(net2987));
 AO21x1_ASAP7_75t_R _08834_ (.A1(_02841_),
    .A2(net5286),
    .B(net5361),
    .Y(_02888_));
 AOI21x1_ASAP7_75t_R _08835_ (.A1(_00258_),
    .A2(net4694),
    .B(_02888_),
    .Y(_00633_));
 AO21x1_ASAP7_75t_R _08836_ (.A1(net4693),
    .A2(_00257_),
    .B(net5361),
    .Y(_02889_));
 AOI21x1_ASAP7_75t_R _08837_ (.A1(net5285),
    .A2(net4631),
    .B(_02889_),
    .Y(_00634_));
 AO21x1_ASAP7_75t_R _08838_ (.A1(net4693),
    .A2(_00256_),
    .B(net5361),
    .Y(_02890_));
 AOI21x1_ASAP7_75t_R _08839_ (.A1(net5284),
    .A2(net4631),
    .B(_02890_),
    .Y(_00635_));
 AO21x1_ASAP7_75t_R _08840_ (.A1(net4695),
    .A2(_00255_),
    .B(net5361),
    .Y(_02891_));
 AOI21x1_ASAP7_75t_R _08841_ (.A1(net5283),
    .A2(net4632),
    .B(_02891_),
    .Y(_00636_));
 AO21x1_ASAP7_75t_R _08842_ (.A1(net4695),
    .A2(_00254_),
    .B(net5361),
    .Y(_02892_));
 AOI21x1_ASAP7_75t_R _08843_ (.A1(net5282),
    .A2(net4632),
    .B(_02892_),
    .Y(_00637_));
 INVx1_ASAP7_75t_R _08844_ (.A(_00365_),
    .Y(_02893_));
 AO21x1_ASAP7_75t_R _08845_ (.A1(net5332),
    .A2(net5329),
    .B(_01124_),
    .Y(_02894_));
 NOR2x1p5_ASAP7_75t_R _08846_ (.A(_02894_),
    .B(_01100_),
    .Y(_02895_));
 INVx2_ASAP7_75t_R _08847_ (.A(_02895_),
    .Y(_02896_));
 OR3x1_ASAP7_75t_R _08848_ (.A(_02896_),
    .B(_01126_),
    .C(_01119_),
    .Y(_02897_));
 BUFx3_ASAP7_75t_R place2986 (.A(_06268_),
    .Y(net2986));
 INVx2_ASAP7_75t_R _08850_ (.A(_02897_),
    .Y(_02899_));
 BUFx3_ASAP7_75t_R place2985 (.A(_06320_),
    .Y(net2985));
 INVx1_ASAP7_75t_R _08852_ (.A(_00482_),
    .Y(_02901_));
 AND3x1_ASAP7_75t_R _08853_ (.A(_02901_),
    .B(net5262),
    .C(net5261),
    .Y(_02902_));
 AO21x1_ASAP7_75t_R _08854_ (.A1(_02902_),
    .A2(net5260),
    .B(net5330),
    .Y(_02903_));
 AO21x1_ASAP7_75t_R _08855_ (.A1(net3998),
    .A2(_02903_),
    .B(net5360),
    .Y(_02904_));
 AO21x1_ASAP7_75t_R _08856_ (.A1(_02893_),
    .A2(net4017),
    .B(_02904_),
    .Y(_00638_));
 INVx1_ASAP7_75t_R _08857_ (.A(_00366_),
    .Y(_02905_));
 NOR2x1_ASAP7_75t_R _08858_ (.A(_00485_),
    .B(\u_fft.sched[42] ),
    .Y(_02906_));
 AND3x1_ASAP7_75t_R _08859_ (.A(net5018),
    .B(net5260),
    .C(net5261),
    .Y(_02907_));
 AO21x1_ASAP7_75t_R _08860_ (.A1(_02906_),
    .A2(net4846),
    .B(net4015),
    .Y(_02908_));
 OA211x2_ASAP7_75t_R _08861_ (.A1(_02905_),
    .A2(net3999),
    .B(_02908_),
    .C(net211),
    .Y(_00639_));
 INVx1_ASAP7_75t_R _08862_ (.A(_00484_),
    .Y(_02909_));
 AND3x1_ASAP7_75t_R _08863_ (.A(net4846),
    .B(_02909_),
    .C(net5262),
    .Y(_02910_));
 OA21x2_ASAP7_75t_R _08864_ (.A1(net5080),
    .A2(net3999),
    .B(net211),
    .Y(_02911_));
 OA21x2_ASAP7_75t_R _08865_ (.A1(net4015),
    .A2(_02910_),
    .B(_02911_),
    .Y(_00640_));
 INVx1_ASAP7_75t_R _08866_ (.A(_02907_),
    .Y(_02912_));
 OAI21x1_ASAP7_75t_R _08867_ (.A1(_00489_),
    .A2(_02912_),
    .B(net3999),
    .Y(_02913_));
 OA211x2_ASAP7_75t_R _08868_ (.A1(net5081),
    .A2(net3999),
    .B(_02913_),
    .C(net211),
    .Y(_00641_));
 BUFx3_ASAP7_75t_R place2984 (.A(net5636),
    .Y(net2984));
 BUFx3_ASAP7_75t_R place2983 (.A(net5894),
    .Y(net2983));
 AND3x1_ASAP7_75t_R _08871_ (.A(_02907_),
    .B(net4847),
    .C(\u_fft.sched[42] ),
    .Y(_02916_));
 OA21x2_ASAP7_75t_R _08872_ (.A1(net4018),
    .A2(_02916_),
    .B(net211),
    .Y(_02917_));
 OA21x2_ASAP7_75t_R _08873_ (.A1(net5079),
    .A2(net3999),
    .B(_02917_),
    .Y(_00642_));
 INVx1_ASAP7_75t_R _08874_ (.A(_00485_),
    .Y(_02918_));
 AND3x1_ASAP7_75t_R _08875_ (.A(_02907_),
    .B(_02918_),
    .C(net5068),
    .Y(_02919_));
 NAND2x1p5_ASAP7_75t_R _08876_ (.A(net5277),
    .B(net4018),
    .Y(_02920_));
 OA211x2_ASAP7_75t_R _08877_ (.A1(net4018),
    .A2(_02919_),
    .B(net211),
    .C(_02920_),
    .Y(_00643_));
 OR3x1_ASAP7_75t_R _08878_ (.A(_02912_),
    .B(_00484_),
    .C(net5262),
    .Y(_02921_));
 AO21x1_ASAP7_75t_R _08879_ (.A1(net5276),
    .A2(net4018),
    .B(net5360),
    .Y(_02922_));
 AOI21x1_ASAP7_75t_R _08880_ (.A1(net6043),
    .A2(_02921_),
    .B(_02922_),
    .Y(_00644_));
 OA21x2_ASAP7_75t_R _08881_ (.A1(_00491_),
    .A2(_02912_),
    .B(net3999),
    .Y(_02923_));
 AOI211x1_ASAP7_75t_R _08882_ (.A1(net5275),
    .A2(net6039),
    .B(_02923_),
    .C(net5360),
    .Y(_00645_));
 INVx1_ASAP7_75t_R _08883_ (.A(net5260),
    .Y(_02924_));
 OR5x1_ASAP7_75t_R _08884_ (.A(_02924_),
    .B(\u_fft.sched[42] ),
    .C(net5330),
    .D(net4869),
    .E(net5261),
    .Y(_02925_));
 AO21x1_ASAP7_75t_R _08885_ (.A1(net5274),
    .A2(net4018),
    .B(net5360),
    .Y(_02926_));
 AOI21x1_ASAP7_75t_R _08886_ (.A1(net6043),
    .A2(_02925_),
    .B(_02926_),
    .Y(_00646_));
 OR5x1_ASAP7_75t_R _08887_ (.A(_02924_),
    .B(\u_fft.sched[42] ),
    .C(net5330),
    .D(_00485_),
    .E(net5261),
    .Y(_02927_));
 AO21x1_ASAP7_75t_R _08888_ (.A1(_00236_),
    .A2(net4018),
    .B(net5360),
    .Y(_02928_));
 AOI21x1_ASAP7_75t_R _08889_ (.A1(net6043),
    .A2(_02927_),
    .B(_02928_),
    .Y(_00647_));
 NOR2x1_ASAP7_75t_R _08890_ (.A(net5262),
    .B(net5261),
    .Y(_02929_));
 NAND2x1_ASAP7_75t_R _08891_ (.A(_00487_),
    .B(_02929_),
    .Y(_02930_));
 XOR2x2_ASAP7_75t_R _08892_ (.A(_02930_),
    .B(net5260),
    .Y(_02931_));
 INVx1_ASAP7_75t_R _08893_ (.A(_02931_),
    .Y(_02932_));
 INVx1_ASAP7_75t_R _08894_ (.A(_00490_),
    .Y(_02933_));
 NOR2x1_ASAP7_75t_R _08895_ (.A(net5260),
    .B(net5263),
    .Y(_02934_));
 AO21x1_ASAP7_75t_R _08896_ (.A1(net4899),
    .A2(_02934_),
    .B(net5264),
    .Y(_02935_));
 INVx1_ASAP7_75t_R _08897_ (.A(_02935_),
    .Y(_02936_));
 AND4x1_ASAP7_75t_R _08898_ (.A(_02932_),
    .B(_00483_),
    .C(_02933_),
    .D(_02936_),
    .Y(_02937_));
 OR3x1_ASAP7_75t_R _08899_ (.A(net5262),
    .B(net5263),
    .C(net5264),
    .Y(_02938_));
 XOR2x2_ASAP7_75t_R _08900_ (.A(_02938_),
    .B(net5261),
    .Y(_02939_));
 INVx1_ASAP7_75t_R _08901_ (.A(_02939_),
    .Y(_02940_));
 AND3x1_ASAP7_75t_R _08902_ (.A(_02937_),
    .B(net5018),
    .C(_02940_),
    .Y(_02941_));
 OA21x2_ASAP7_75t_R _08903_ (.A1(net4016),
    .A2(_02941_),
    .B(net211),
    .Y(_02942_));
 OA21x2_ASAP7_75t_R _08904_ (.A1(net5070),
    .A2(net6035),
    .B(_02942_),
    .Y(_00648_));
 AND3x1_ASAP7_75t_R _08905_ (.A(_02932_),
    .B(_02901_),
    .C(_02933_),
    .Y(_02943_));
 AO21x1_ASAP7_75t_R _08906_ (.A1(_02943_),
    .A2(_02940_),
    .B(net5330),
    .Y(_02944_));
 AO21x1_ASAP7_75t_R _08907_ (.A1(net3998),
    .A2(_02944_),
    .B(net5360),
    .Y(_02945_));
 AO21x1_ASAP7_75t_R _08908_ (.A1(net5071),
    .A2(net4016),
    .B(_02945_),
    .Y(_00649_));
 OR3x1_ASAP7_75t_R _08909_ (.A(_02931_),
    .B(net5330),
    .C(net4643),
    .Y(_02946_));
 INVx1_ASAP7_75t_R _08910_ (.A(_00483_),
    .Y(_02947_));
 NAND2x1_ASAP7_75t_R _08911_ (.A(_02947_),
    .B(net4735),
    .Y(_02948_));
 OR3x1_ASAP7_75t_R _08912_ (.A(_02946_),
    .B(net4844),
    .C(_02948_),
    .Y(_02949_));
 AO21x1_ASAP7_75t_R _08913_ (.A1(net5272),
    .A2(net4016),
    .B(net5360),
    .Y(_02950_));
 AOI21x1_ASAP7_75t_R _08914_ (.A1(net6036),
    .A2(_02949_),
    .B(_02950_),
    .Y(_00650_));
 OR3x1_ASAP7_75t_R _08915_ (.A(_02946_),
    .B(_00484_),
    .C(net4844),
    .Y(_02951_));
 AO21x1_ASAP7_75t_R _08916_ (.A1(net5271),
    .A2(net4016),
    .B(net5360),
    .Y(_02952_));
 AOI21x1_ASAP7_75t_R _08917_ (.A1(net6033),
    .A2(_02951_),
    .B(_02952_),
    .Y(_00651_));
 OR3x1_ASAP7_75t_R _08918_ (.A(_02931_),
    .B(net5330),
    .C(_02933_),
    .Y(_02953_));
 OR4x1_ASAP7_75t_R _08919_ (.A(_02953_),
    .B(_02947_),
    .C(_02939_),
    .D(net4845),
    .Y(_02954_));
 BUFx3_ASAP7_75t_R place2982 (.A(_02244_),
    .Y(net2982));
 AO21x1_ASAP7_75t_R _08921_ (.A1(net3998),
    .A2(_02954_),
    .B(net5360),
    .Y(_02956_));
 AOI21x1_ASAP7_75t_R _08922_ (.A1(net6028),
    .A2(net5270),
    .B(_02956_),
    .Y(_00652_));
 OR3x1_ASAP7_75t_R _08923_ (.A(_02953_),
    .B(net4869),
    .C(net4844),
    .Y(_02957_));
 AO21x1_ASAP7_75t_R _08924_ (.A1(net5269),
    .A2(net4016),
    .B(net5360),
    .Y(_02958_));
 AOI21x1_ASAP7_75t_R _08925_ (.A1(net6037),
    .A2(_02957_),
    .B(_02958_),
    .Y(_00653_));
 OR3x1_ASAP7_75t_R _08926_ (.A(_02953_),
    .B(net4843),
    .C(_02948_),
    .Y(_02959_));
 AO21x1_ASAP7_75t_R _08927_ (.A1(net6037),
    .A2(_02959_),
    .B(net5360),
    .Y(_02960_));
 AOI21x1_ASAP7_75t_R _08928_ (.A1(net5268),
    .A2(net6028),
    .B(_02960_),
    .Y(_00654_));
 OR3x1_ASAP7_75t_R _08929_ (.A(_02953_),
    .B(_00484_),
    .C(net4843),
    .Y(_02961_));
 AO21x1_ASAP7_75t_R _08930_ (.A1(net5267),
    .A2(net4016),
    .B(net5360),
    .Y(_02962_));
 AOI21x1_ASAP7_75t_R _08931_ (.A1(net6034),
    .A2(_02961_),
    .B(_02962_),
    .Y(_00655_));
 AND3x4_ASAP7_75t_R _08932_ (.A(_02899_),
    .B(net5018),
    .C(_02939_),
    .Y(_02963_));
 NOR2x1_ASAP7_75t_R _08933_ (.A(net5266),
    .B(net3998),
    .Y(_02964_));
 AO21x1_ASAP7_75t_R _08934_ (.A1(_02963_),
    .A2(net4527),
    .B(_02964_),
    .Y(_02965_));
 AND2x2_ASAP7_75t_R _08935_ (.A(_02965_),
    .B(net211),
    .Y(_00656_));
 NOR2x1_ASAP7_75t_R _08936_ (.A(net5265),
    .B(net3998),
    .Y(_02966_));
 AO21x1_ASAP7_75t_R _08937_ (.A1(_02963_),
    .A2(_02943_),
    .B(_02966_),
    .Y(_02967_));
 AND2x2_ASAP7_75t_R _08938_ (.A(_02967_),
    .B(net211),
    .Y(_00657_));
 NAND2x1_ASAP7_75t_R _08939_ (.A(net5018),
    .B(net5066),
    .Y(_02968_));
 AO21x1_ASAP7_75t_R _08940_ (.A1(net5066),
    .A2(net4017),
    .B(net5360),
    .Y(_02969_));
 AO21x1_ASAP7_75t_R _08941_ (.A1(net6037),
    .A2(_02968_),
    .B(_02969_),
    .Y(_00658_));
 AND3x1_ASAP7_75t_R _08942_ (.A(_02947_),
    .B(net5018),
    .C(_02899_),
    .Y(_02970_));
 AO21x1_ASAP7_75t_R _08943_ (.A1(net5067),
    .A2(net4015),
    .B(_02970_),
    .Y(_02971_));
 AND2x2_ASAP7_75t_R _08944_ (.A(_02971_),
    .B(net211),
    .Y(_00659_));
 AND3x1_ASAP7_75t_R _08945_ (.A(net4643),
    .B(net5018),
    .C(_02899_),
    .Y(_02972_));
 AO21x1_ASAP7_75t_R _08946_ (.A1(net5069),
    .A2(net4017),
    .B(_02972_),
    .Y(_02973_));
 AND2x2_ASAP7_75t_R _08947_ (.A(_02973_),
    .B(net5363),
    .Y(_00660_));
 NOR2x1_ASAP7_75t_R _08948_ (.A(net5261),
    .B(net3998),
    .Y(_02974_));
 OA21x2_ASAP7_75t_R _08949_ (.A1(_02974_),
    .A2(_02963_),
    .B(net211),
    .Y(_00661_));
 AND3x1_ASAP7_75t_R _08950_ (.A(net4017),
    .B(net5363),
    .C(net4900),
    .Y(_00662_));
 NOR2x2_ASAP7_75t_R _08951_ (.A(net5360),
    .B(net4085),
    .Y(_02975_));
 NAND2x1_ASAP7_75t_R _08952_ (.A(net5258),
    .B(net4737),
    .Y(_02976_));
 INVx1_ASAP7_75t_R _08953_ (.A(net4736),
    .Y(_02977_));
 NAND2x1_ASAP7_75t_R _08954_ (.A(\u_fft.sched[45] ),
    .B(net4683),
    .Y(_02978_));
 AND3x1_ASAP7_75t_R _08955_ (.A(net4042),
    .B(_02976_),
    .C(_02978_),
    .Y(_00663_));
 INVx1_ASAP7_75t_R _08956_ (.A(_00493_),
    .Y(_02979_));
 AND3x1_ASAP7_75t_R _08957_ (.A(net4152),
    .B(_02979_),
    .C(net4683),
    .Y(_02980_));
 NOR2x1_ASAP7_75t_R _08958_ (.A(net5257),
    .B(net4683),
    .Y(_02981_));
 OA21x2_ASAP7_75t_R _08959_ (.A1(_02980_),
    .A2(_02981_),
    .B(net211),
    .Y(_00664_));
 INVx1_ASAP7_75t_R _08960_ (.A(_00492_),
    .Y(_02982_));
 AND3x1_ASAP7_75t_R _08961_ (.A(_02977_),
    .B(net5000),
    .C(_02982_),
    .Y(_02983_));
 INVx1_ASAP7_75t_R _08962_ (.A(_02983_),
    .Y(_02984_));
 AO21x1_ASAP7_75t_R _08963_ (.A1(net4683),
    .A2(_02982_),
    .B(net5000),
    .Y(_02985_));
 AND3x1_ASAP7_75t_R _08964_ (.A(net4042),
    .B(net4572),
    .C(_02985_),
    .Y(_00665_));
 AND3x1_ASAP7_75t_R _08965_ (.A(net5000),
    .B(net4999),
    .C(\u_fft.sched[45] ),
    .Y(_02986_));
 INVx1_ASAP7_75t_R _08966_ (.A(_02986_),
    .Y(_02987_));
 OR3x1_ASAP7_75t_R _08967_ (.A(net4737),
    .B(net5256),
    .C(_02987_),
    .Y(_02988_));
 AO21x1_ASAP7_75t_R _08968_ (.A1(net4682),
    .A2(_02986_),
    .B(net4998),
    .Y(_02989_));
 AND3x1_ASAP7_75t_R _08969_ (.A(net4042),
    .B(_02988_),
    .C(_02989_),
    .Y(_00666_));
 NOR2x1_ASAP7_75t_R _08970_ (.A(net5255),
    .B(net5256),
    .Y(_02990_));
 INVx1_ASAP7_75t_R _08971_ (.A(net4897),
    .Y(_02991_));
 AO21x1_ASAP7_75t_R _08972_ (.A1(net4629),
    .A2(net4998),
    .B(\u_fft.sched[49] ),
    .Y(_02992_));
 OA211x2_ASAP7_75t_R _08973_ (.A1(net4572),
    .A2(_02991_),
    .B(_02975_),
    .C(_02992_),
    .Y(_00667_));
 NAND2x1_ASAP7_75t_R _08974_ (.A(\u_fft.sched[50] ),
    .B(net4898),
    .Y(_02993_));
 OA211x2_ASAP7_75t_R _08975_ (.A1(_02987_),
    .A2(net4842),
    .B(net4152),
    .C(net4683),
    .Y(_02994_));
 NOR2x1_ASAP7_75t_R _08976_ (.A(_00064_),
    .B(net4683),
    .Y(_02995_));
 AO21x1_ASAP7_75t_R _08977_ (.A1(_02986_),
    .A2(net4897),
    .B(\u_fft.sched[50] ),
    .Y(_02996_));
 OA211x2_ASAP7_75t_R _08978_ (.A1(_02994_),
    .A2(_02995_),
    .B(net211),
    .C(_02996_),
    .Y(_00668_));
 NOR2x1_ASAP7_75t_R _08979_ (.A(_02993_),
    .B(_02984_),
    .Y(_02997_));
 XOR2x2_ASAP7_75t_R _08980_ (.A(net4526),
    .B(net5254),
    .Y(_02998_));
 INVx3_ASAP7_75t_R _08981_ (.A(_02975_),
    .Y(_02999_));
 NOR2x1_ASAP7_75t_R _08982_ (.A(_02998_),
    .B(_02999_),
    .Y(_00669_));
 AND5x1_ASAP7_75t_R _08983_ (.A(\u_fft.sched[50] ),
    .B(net4682),
    .C(net4997),
    .D(_02986_),
    .E(_02990_),
    .Y(_03000_));
 XOR2x2_ASAP7_75t_R _08984_ (.A(net4628),
    .B(net5253),
    .Y(_03001_));
 NOR2x1_ASAP7_75t_R _08985_ (.A(_03001_),
    .B(_02999_),
    .Y(_00670_));
 AND3x1_ASAP7_75t_R _08986_ (.A(_02997_),
    .B(net4997),
    .C(net4996),
    .Y(_03002_));
 XOR2x2_ASAP7_75t_R _08987_ (.A(_03002_),
    .B(net5252),
    .Y(_03003_));
 NOR2x1_ASAP7_75t_R _08988_ (.A(_03003_),
    .B(_02999_),
    .Y(_00671_));
 AND3x1_ASAP7_75t_R _08989_ (.A(_03000_),
    .B(\u_fft.sched[53] ),
    .C(net4996),
    .Y(_03004_));
 XOR2x2_ASAP7_75t_R _08990_ (.A(_03004_),
    .B(net5251),
    .Y(_03005_));
 NOR2x1_ASAP7_75t_R _08991_ (.A(_03005_),
    .B(_02999_),
    .Y(_00672_));
 BUFx3_ASAP7_75t_R place2981 (.A(_02261_),
    .Y(net2981));
 AND2x2_ASAP7_75t_R _08993_ (.A(net211),
    .B(_00496_),
    .Y(_03007_));
 AO32x1_ASAP7_75t_R _08994_ (.A1(net4179),
    .A2(net4086),
    .A3(_03007_),
    .B1(\u_fft.sched[55] ),
    .B2(_02975_),
    .Y(_00673_));
 NOR2x1_ASAP7_75t_R _08995_ (.A(_00340_),
    .B(net5360),
    .Y(_03008_));
 AO32x1_ASAP7_75t_R _08996_ (.A1(net4179),
    .A2(net4086),
    .A3(_03008_),
    .B1(_02975_),
    .B2(net4927),
    .Y(_00674_));
 XOR2x2_ASAP7_75t_R _08997_ (.A(net4659),
    .B(net4758),
    .Y(_03009_));
 AO21x1_ASAP7_75t_R _08998_ (.A1(net4179),
    .A2(_03009_),
    .B(net4043),
    .Y(_03010_));
 BUFx3_ASAP7_75t_R place2980 (.A(_03965_),
    .Y(net2980));
 OA211x2_ASAP7_75t_R _09000_ (.A1(\u_fft.sched[57] ),
    .A2(net4086),
    .B(_03010_),
    .C(net5362),
    .Y(_00675_));
 OAI21x1_ASAP7_75t_R _09001_ (.A1(net4757),
    .A2(_00498_),
    .B(_00500_),
    .Y(_03012_));
 INVx1_ASAP7_75t_R _09002_ (.A(_00501_),
    .Y(_03013_));
 INVx1_ASAP7_75t_R _09003_ (.A(_00499_),
    .Y(_03014_));
 AND3x1_ASAP7_75t_R _09004_ (.A(_03013_),
    .B(_03014_),
    .C(_00338_),
    .Y(_03015_));
 NOR2x1_ASAP7_75t_R _09005_ (.A(_03012_),
    .B(_03015_),
    .Y(_03016_));
 XOR2x2_ASAP7_75t_R _09006_ (.A(net4578),
    .B(net4756),
    .Y(_03017_));
 AO21x1_ASAP7_75t_R _09007_ (.A1(net4179),
    .A2(_03017_),
    .B(net4043),
    .Y(_03018_));
 OA211x2_ASAP7_75t_R _09008_ (.A1(net4086),
    .A2(net4928),
    .B(_03018_),
    .C(net5362),
    .Y(_00676_));
 OA21x2_ASAP7_75t_R _09009_ (.A1(_00339_),
    .A2(net4758),
    .B(_00500_),
    .Y(_03019_));
 OAI21x1_ASAP7_75t_R _09010_ (.A1(_00503_),
    .A2(_03019_),
    .B(_00502_),
    .Y(_03020_));
 INVx1_ASAP7_75t_R _09011_ (.A(_00505_),
    .Y(_03021_));
 XOR2x2_ASAP7_75t_R _09012_ (.A(net4571),
    .B(net4705),
    .Y(_03022_));
 AO21x1_ASAP7_75t_R _09013_ (.A1(net4179),
    .A2(_03022_),
    .B(net4043),
    .Y(_03023_));
 OA211x2_ASAP7_75t_R _09014_ (.A1(net4086),
    .A2(net4929),
    .B(_03023_),
    .C(net5362),
    .Y(_00677_));
 OAI21x1_ASAP7_75t_R _09015_ (.A1(_00503_),
    .A2(_03016_),
    .B(_00502_),
    .Y(_03024_));
 INVx1_ASAP7_75t_R _09016_ (.A(_00504_),
    .Y(_03025_));
 AO21x1_ASAP7_75t_R _09017_ (.A1(_03024_),
    .A2(_03021_),
    .B(_03025_),
    .Y(_03026_));
 INVx1_ASAP7_75t_R _09018_ (.A(_00507_),
    .Y(_03027_));
 XOR2x2_ASAP7_75t_R _09019_ (.A(net4473),
    .B(net4704),
    .Y(_03028_));
 AO21x1_ASAP7_75t_R _09020_ (.A1(net4179),
    .A2(_03028_),
    .B(net4043),
    .Y(_03029_));
 OA211x2_ASAP7_75t_R _09021_ (.A1(net4930),
    .A2(net4086),
    .B(_03029_),
    .C(net5362),
    .Y(_00678_));
 AO21x1_ASAP7_75t_R _09022_ (.A1(_03020_),
    .A2(_03021_),
    .B(_03025_),
    .Y(_03030_));
 INVx1_ASAP7_75t_R _09023_ (.A(_00506_),
    .Y(_03031_));
 AO21x1_ASAP7_75t_R _09024_ (.A1(_03030_),
    .A2(_03027_),
    .B(_03031_),
    .Y(_03032_));
 INVx1_ASAP7_75t_R _09025_ (.A(_00509_),
    .Y(_03033_));
 XOR2x2_ASAP7_75t_R _09026_ (.A(net4470),
    .B(net4703),
    .Y(_03034_));
 AO21x1_ASAP7_75t_R _09027_ (.A1(net4179),
    .A2(_03034_),
    .B(net4043),
    .Y(_03035_));
 OA211x2_ASAP7_75t_R _09028_ (.A1(net4931),
    .A2(net4086),
    .B(_03035_),
    .C(net5362),
    .Y(_00679_));
 AO21x1_ASAP7_75t_R _09029_ (.A1(_03026_),
    .A2(_03027_),
    .B(_03031_),
    .Y(_03036_));
 INVx1_ASAP7_75t_R _09030_ (.A(_00508_),
    .Y(_03037_));
 AO21x1_ASAP7_75t_R _09031_ (.A1(_03036_),
    .A2(_03033_),
    .B(_03037_),
    .Y(_03038_));
 INVx1_ASAP7_75t_R _09032_ (.A(_00511_),
    .Y(_03039_));
 XOR2x2_ASAP7_75t_R _09033_ (.A(net4375),
    .B(net4702),
    .Y(_03040_));
 AO21x1_ASAP7_75t_R _09034_ (.A1(net4179),
    .A2(_03040_),
    .B(net4043),
    .Y(_03041_));
 OA211x2_ASAP7_75t_R _09035_ (.A1(\u_fft.sched[62] ),
    .A2(net4086),
    .B(_03041_),
    .C(net5362),
    .Y(_00680_));
 AO21x1_ASAP7_75t_R _09036_ (.A1(_03032_),
    .A2(_03033_),
    .B(_03037_),
    .Y(_03042_));
 INVx1_ASAP7_75t_R _09037_ (.A(_00510_),
    .Y(_03043_));
 AO21x1_ASAP7_75t_R _09038_ (.A1(_03042_),
    .A2(_03039_),
    .B(_03043_),
    .Y(_03044_));
 XNOR2x2_ASAP7_75t_R _09039_ (.A(net4755),
    .B(_03044_),
    .Y(_03045_));
 AO21x1_ASAP7_75t_R _09040_ (.A1(net4179),
    .A2(_03045_),
    .B(net4043),
    .Y(_03046_));
 OA211x2_ASAP7_75t_R _09041_ (.A1(net4932),
    .A2(net4086),
    .B(_03046_),
    .C(net5362),
    .Y(_00681_));
 NAND2x1_ASAP7_75t_R _09042_ (.A(_03039_),
    .B(_03038_),
    .Y(_03047_));
 AO21x1_ASAP7_75t_R _09043_ (.A1(_03047_),
    .A2(_00510_),
    .B(_00513_),
    .Y(_03048_));
 NAND2x1_ASAP7_75t_R _09044_ (.A(_00512_),
    .B(_03048_),
    .Y(_03049_));
 XOR2x2_ASAP7_75t_R _09045_ (.A(net5250),
    .B(net5265),
    .Y(_03050_));
 OAI21x1_ASAP7_75t_R _09046_ (.A1(_03050_),
    .A2(_03049_),
    .B(net211),
    .Y(_03051_));
 AOI21x1_ASAP7_75t_R _09047_ (.A1(_03049_),
    .A2(_03050_),
    .B(_03051_),
    .Y(_03052_));
 AO32x1_ASAP7_75t_R _09048_ (.A1(net4179),
    .A2(net4086),
    .A3(_03052_),
    .B1(_02975_),
    .B2(\u_fft.sched[64] ),
    .Y(_00682_));
 NOR2x1_ASAP7_75t_R _09049_ (.A(net5360),
    .B(_00176_),
    .Y(_00715_));
 AND2x2_ASAP7_75t_R _09050_ (.A(_00046_),
    .B(_00328_),
    .Y(_03053_));
 BUFx3_ASAP7_75t_R place2979 (.A(_03975_),
    .Y(net2979));
 INVx1_ASAP7_75t_R _09052_ (.A(_03053_),
    .Y(_03055_));
 AO21x1_ASAP7_75t_R _09053_ (.A1(_03055_),
    .A2(net5213),
    .B(_00930_),
    .Y(_03056_));
 AND2x2_ASAP7_75t_R _09054_ (.A(_02513_),
    .B(_03056_),
    .Y(_03057_));
 BUFx3_ASAP7_75t_R place2978 (.A(_03983_),
    .Y(net2978));
 INVx1_ASAP7_75t_R _09056_ (.A(_03057_),
    .Y(_03059_));
 INVx1_ASAP7_75t_R _09057_ (.A(net2725),
    .Y(_03060_));
 INVx1_ASAP7_75t_R _09058_ (.A(_02443_),
    .Y(_03061_));
 NAND2x1_ASAP7_75t_R _09059_ (.A(_02452_),
    .B(_02413_),
    .Y(_03062_));
 NOR2x1_ASAP7_75t_R _09060_ (.A(_03061_),
    .B(_03062_),
    .Y(_03063_));
 AOI21x1_ASAP7_75t_R _09061_ (.A1(_03060_),
    .A2(_03063_),
    .B(net5144),
    .Y(_03064_));
 AOI21x1_ASAP7_75t_R _09062_ (.A1(net4642),
    .A2(_03064_),
    .B(_00046_),
    .Y(_03065_));
 OAI21x1_ASAP7_75t_R _09063_ (.A1(net4570),
    .A2(net2703),
    .B(net4995),
    .Y(_03066_));
 NOR2x1_ASAP7_75t_R _09064_ (.A(net4995),
    .B(net4896),
    .Y(_03067_));
 NAND3x2_ASAP7_75t_R _09065_ (.B(net4626),
    .C(_03067_),
    .Y(_03068_),
    .A(net2711));
 AOI21x1_ASAP7_75t_R _09066_ (.A1(_03066_),
    .A2(_03068_),
    .B(net5360),
    .Y(_00716_));
 OAI21x1_ASAP7_75t_R _09067_ (.A1(net4570),
    .A2(net2703),
    .B(net5044),
    .Y(_03069_));
 NOR2x1_ASAP7_75t_R _09068_ (.A(_00517_),
    .B(net4896),
    .Y(_03070_));
 NAND3x2_ASAP7_75t_R _09069_ (.B(net4626),
    .C(_03070_),
    .Y(_03071_),
    .A(net5418));
 AOI21x1_ASAP7_75t_R _09070_ (.A1(_03069_),
    .A2(_03071_),
    .B(net5360),
    .Y(_00717_));
 INVx1_ASAP7_75t_R _09071_ (.A(net5219),
    .Y(_03072_));
 OAI21x1_ASAP7_75t_R _09072_ (.A1(net4570),
    .A2(net2703),
    .B(_03072_),
    .Y(_03073_));
 XNOR2x2_ASAP7_75t_R _09073_ (.A(net5219),
    .B(net4820),
    .Y(_03074_));
 NOR2x1_ASAP7_75t_R _09074_ (.A(net4896),
    .B(_03074_),
    .Y(_03075_));
 NAND3x2_ASAP7_75t_R _09075_ (.B(net4625),
    .C(_03075_),
    .Y(_03076_),
    .A(net2711));
 AOI21x1_ASAP7_75t_R _09076_ (.A1(_03073_),
    .A2(_03076_),
    .B(net5360),
    .Y(_00718_));
 INVx1_ASAP7_75t_R _09077_ (.A(net5218),
    .Y(_03077_));
 OAI21x1_ASAP7_75t_R _09078_ (.A1(net4570),
    .A2(net2703),
    .B(net4895),
    .Y(_03078_));
 OR3x1_ASAP7_75t_R _09079_ (.A(net5221),
    .B(net5219),
    .C(net5220),
    .Y(_03079_));
 XOR2x2_ASAP7_75t_R _09080_ (.A(_03079_),
    .B(_03077_),
    .Y(_03080_));
 NOR2x1_ASAP7_75t_R _09081_ (.A(net4896),
    .B(_03080_),
    .Y(_03081_));
 NAND3x2_ASAP7_75t_R _09082_ (.B(net5418),
    .C(_03081_),
    .Y(_03082_),
    .A(net4625));
 AOI21x1_ASAP7_75t_R _09083_ (.A1(_03078_),
    .A2(_03082_),
    .B(net5360),
    .Y(_00719_));
 INVx1_ASAP7_75t_R _09084_ (.A(_00180_),
    .Y(_03083_));
 OAI21x1_ASAP7_75t_R _09085_ (.A1(net4570),
    .A2(net2703),
    .B(net4894),
    .Y(_03084_));
 OR3x1_ASAP7_75t_R _09086_ (.A(net5218),
    .B(net5219),
    .C(net4820),
    .Y(_03085_));
 XOR2x2_ASAP7_75t_R _09087_ (.A(_03085_),
    .B(_03083_),
    .Y(_03086_));
 NOR2x1_ASAP7_75t_R _09088_ (.A(net4896),
    .B(_03086_),
    .Y(_03087_));
 NAND3x1_ASAP7_75t_R _09089_ (.A(net5418),
    .B(net4625),
    .C(_03087_),
    .Y(_03088_));
 AOI21x1_ASAP7_75t_R _09090_ (.A1(_03084_),
    .A2(_03088_),
    .B(net5360),
    .Y(_00720_));
 INVx1_ASAP7_75t_R _09091_ (.A(net5217),
    .Y(_03089_));
 OAI21x1_ASAP7_75t_R _09092_ (.A1(net4569),
    .A2(net2703),
    .B(net4893),
    .Y(_03090_));
 XOR2x2_ASAP7_75t_R _09093_ (.A(net4860),
    .B(_03089_),
    .Y(_03091_));
 NOR2x1_ASAP7_75t_R _09094_ (.A(net4896),
    .B(_03091_),
    .Y(_03092_));
 NAND3x2_ASAP7_75t_R _09095_ (.B(net4626),
    .C(_03092_),
    .Y(_03093_),
    .A(net2711));
 AOI21x1_ASAP7_75t_R _09096_ (.A1(_03090_),
    .A2(_03093_),
    .B(net5360),
    .Y(_00721_));
 INVx1_ASAP7_75t_R _09097_ (.A(net5216),
    .Y(_03094_));
 OAI21x1_ASAP7_75t_R _09098_ (.A1(net4569),
    .A2(net2703),
    .B(net4892),
    .Y(_03095_));
 OR3x1_ASAP7_75t_R _09099_ (.A(net5043),
    .B(net5217),
    .C(_00516_),
    .Y(_03096_));
 XOR2x2_ASAP7_75t_R _09100_ (.A(net4734),
    .B(_03094_),
    .Y(_03097_));
 NOR2x1_ASAP7_75t_R _09101_ (.A(net4896),
    .B(_03097_),
    .Y(_03098_));
 NAND3x1_ASAP7_75t_R _09102_ (.A(net5418),
    .B(net4626),
    .C(_03098_),
    .Y(_03099_));
 AOI21x1_ASAP7_75t_R _09103_ (.A1(_03095_),
    .A2(_03099_),
    .B(net5360),
    .Y(_00722_));
 INVx1_ASAP7_75t_R _09104_ (.A(net5215),
    .Y(_03100_));
 OAI21x1_ASAP7_75t_R _09105_ (.A1(net4570),
    .A2(net2703),
    .B(net4891),
    .Y(_03101_));
 XOR2x2_ASAP7_75t_R _09106_ (.A(net4750),
    .B(_03100_),
    .Y(_03102_));
 NOR2x1_ASAP7_75t_R _09107_ (.A(net4896),
    .B(_03102_),
    .Y(_03103_));
 NAND3x2_ASAP7_75t_R _09108_ (.B(net4627),
    .C(_03103_),
    .Y(_03104_),
    .A(net2711));
 AOI21x1_ASAP7_75t_R _09109_ (.A1(_03101_),
    .A2(_03104_),
    .B(net5360),
    .Y(_00723_));
 INVx1_ASAP7_75t_R _09110_ (.A(net5214),
    .Y(_03105_));
 OAI21x1_ASAP7_75t_R _09111_ (.A1(net4570),
    .A2(net2703),
    .B(net4890),
    .Y(_03106_));
 OR3x1_ASAP7_75t_R _09112_ (.A(_03096_),
    .B(net5215),
    .C(net5216),
    .Y(_03107_));
 XOR2x2_ASAP7_75t_R _09113_ (.A(_03107_),
    .B(_03105_),
    .Y(_03108_));
 NOR2x1_ASAP7_75t_R _09114_ (.A(net4896),
    .B(_03108_),
    .Y(_03109_));
 NAND3x2_ASAP7_75t_R _09115_ (.B(net4627),
    .C(_03109_),
    .Y(_03110_),
    .A(net2711));
 BUFx3_ASAP7_75t_R place2989 (.A(_05182_),
    .Y(net2989));
 BUFx3_ASAP7_75t_R place2976 (.A(_05151_),
    .Y(net2976));
 AOI21x1_ASAP7_75t_R _09118_ (.A1(_03106_),
    .A2(_03110_),
    .B(net5360),
    .Y(_00724_));
 AND2x2_ASAP7_75t_R _09119_ (.A(_00931_),
    .B(net5363),
    .Y(_00725_));
 AND2x2_ASAP7_75t_R _09120_ (.A(_00331_),
    .B(_00332_),
    .Y(_03113_));
 AO21x1_ASAP7_75t_R _09121_ (.A1(_00898_),
    .A2(_00894_),
    .B(_03113_),
    .Y(_03114_));
 AO21x1_ASAP7_75t_R _09122_ (.A1(_02517_),
    .A2(_00911_),
    .B(_03114_),
    .Y(_03115_));
 INVx2_ASAP7_75t_R _09123_ (.A(_03115_),
    .Y(_03116_));
 OA21x2_ASAP7_75t_R _09124_ (.A1(net4681),
    .A2(\u_mel.k_next[0] ),
    .B(net5362),
    .Y(_03117_));
 OA21x2_ASAP7_75t_R _09125_ (.A1(\u_mel.k[0] ),
    .A2(net4624),
    .B(_03117_),
    .Y(_00726_));
 AO21x1_ASAP7_75t_R _09126_ (.A1(net5211),
    .A2(net4681),
    .B(net5361),
    .Y(_03118_));
 AOI21x1_ASAP7_75t_R _09127_ (.A1(_00555_),
    .A2(net4624),
    .B(_03118_),
    .Y(_00727_));
 INVx1_ASAP7_75t_R _09128_ (.A(_00556_),
    .Y(_03119_));
 AND3x1_ASAP7_75t_R _09129_ (.A(_03119_),
    .B(net5058),
    .C(_03116_),
    .Y(_03120_));
 INVx1_ASAP7_75t_R _09130_ (.A(net4568),
    .Y(_03121_));
 AO21x1_ASAP7_75t_R _09131_ (.A1(net4624),
    .A2(_03119_),
    .B(net5058),
    .Y(_03122_));
 AND3x1_ASAP7_75t_R _09132_ (.A(_03121_),
    .B(net5362),
    .C(_03122_),
    .Y(_00728_));
 AND3x1_ASAP7_75t_R _09133_ (.A(net5058),
    .B(\u_mel.k[1] ),
    .C(\u_mel.k[0] ),
    .Y(_03123_));
 AND2x2_ASAP7_75t_R _09134_ (.A(net4624),
    .B(_03123_),
    .Y(_03124_));
 AND3x4_ASAP7_75t_R _09135_ (.A(net4624),
    .B(net5059),
    .C(_03123_),
    .Y(_03125_));
 NOR2x1p5_ASAP7_75t_R _09136_ (.A(net5361),
    .B(net4567),
    .Y(_03126_));
 OA21x2_ASAP7_75t_R _09137_ (.A1(net5059),
    .A2(_03124_),
    .B(_03126_),
    .Y(_00729_));
 AND3x1_ASAP7_75t_R _09138_ (.A(_03120_),
    .B(net5060),
    .C(net5059),
    .Y(_03127_));
 INVx1_ASAP7_75t_R _09139_ (.A(net4525),
    .Y(_03128_));
 AO21x1_ASAP7_75t_R _09140_ (.A1(net4568),
    .A2(net5059),
    .B(net5060),
    .Y(_03129_));
 AND3x1_ASAP7_75t_R _09141_ (.A(_03128_),
    .B(net5362),
    .C(_03129_),
    .Y(_00730_));
 AND3x1_ASAP7_75t_R _09142_ (.A(_03125_),
    .B(net5062),
    .C(net5060),
    .Y(_03130_));
 INVx1_ASAP7_75t_R _09143_ (.A(_03130_),
    .Y(_03131_));
 AO21x1_ASAP7_75t_R _09144_ (.A1(net4567),
    .A2(net5060),
    .B(net5062),
    .Y(_03132_));
 AND3x1_ASAP7_75t_R _09145_ (.A(_03131_),
    .B(net5362),
    .C(_03132_),
    .Y(_00731_));
 AND3x1_ASAP7_75t_R _09146_ (.A(_03127_),
    .B(net5061),
    .C(net5062),
    .Y(_03133_));
 INVx1_ASAP7_75t_R _09147_ (.A(_03133_),
    .Y(_03134_));
 AO21x1_ASAP7_75t_R _09148_ (.A1(net4525),
    .A2(net5062),
    .B(net5061),
    .Y(_03135_));
 AND3x1_ASAP7_75t_R _09149_ (.A(net4429),
    .B(net5362),
    .C(_03135_),
    .Y(_00732_));
 OR3x1_ASAP7_75t_R _09150_ (.A(_03131_),
    .B(net5210),
    .C(_00170_),
    .Y(_03136_));
 AO21x1_ASAP7_75t_R _09151_ (.A1(_03130_),
    .A2(net5061),
    .B(_00905_),
    .Y(_03137_));
 AND3x1_ASAP7_75t_R _09152_ (.A(_03136_),
    .B(net5362),
    .C(_03137_),
    .Y(_00733_));
 OR3x1_ASAP7_75t_R _09153_ (.A(_03134_),
    .B(_00168_),
    .C(net5210),
    .Y(_03138_));
 AO21x1_ASAP7_75t_R _09154_ (.A1(_03133_),
    .A2(_00905_),
    .B(_00904_),
    .Y(_03139_));
 AND3x1_ASAP7_75t_R _09155_ (.A(_03138_),
    .B(net5362),
    .C(_03139_),
    .Y(_00734_));
 NOR2x1_ASAP7_75t_R _09156_ (.A(net5361),
    .B(net4862),
    .Y(_00735_));
 AND2x2_ASAP7_75t_R _09157_ (.A(net5204),
    .B(_00330_),
    .Y(_03140_));
 INVx2_ASAP7_75t_R _09158_ (.A(_00163_),
    .Y(_03141_));
 OA21x2_ASAP7_75t_R _09159_ (.A1(\mel_ptr[0] ),
    .A2(net4889),
    .B(net5362),
    .Y(_03142_));
 OA21x2_ASAP7_75t_R _09160_ (.A1(_00518_),
    .A2(_03140_),
    .B(_03142_),
    .Y(_00736_));
 INVx1_ASAP7_75t_R _09161_ (.A(_00521_),
    .Y(_03143_));
 AO22x1_ASAP7_75t_R _09162_ (.A1(_03143_),
    .A2(net4889),
    .B1(_03140_),
    .B2(\mel_ptr[1] ),
    .Y(_03144_));
 AND2x2_ASAP7_75t_R _09163_ (.A(_03144_),
    .B(net5362),
    .Y(_00737_));
 NOR2x1_ASAP7_75t_R _09164_ (.A(net5209),
    .B(_00522_),
    .Y(_03145_));
 NAND2x1_ASAP7_75t_R _09165_ (.A(_00900_),
    .B(_03140_),
    .Y(_03146_));
 OA21x2_ASAP7_75t_R _09166_ (.A1(net5204),
    .A2(_03145_),
    .B(_03146_),
    .Y(_03147_));
 AOI211x1_ASAP7_75t_R _09167_ (.A1(net5209),
    .A2(net4819),
    .B(_03147_),
    .C(net5361),
    .Y(_00738_));
 AND4x1_ASAP7_75t_R _09168_ (.A(_03141_),
    .B(_00900_),
    .C(\mel_ptr[1] ),
    .D(\mel_ptr[0] ),
    .Y(_03148_));
 NOR2x1_ASAP7_75t_R _09169_ (.A(_00330_),
    .B(net4889),
    .Y(_03149_));
 NOR2x1_ASAP7_75t_R _09170_ (.A(net5208),
    .B(_03149_),
    .Y(_03150_));
 NAND2x1_ASAP7_75t_R _09171_ (.A(_03148_),
    .B(net5063),
    .Y(_03151_));
 OA211x2_ASAP7_75t_R _09172_ (.A1(_03148_),
    .A2(_03150_),
    .B(_03151_),
    .C(net5362),
    .Y(_00739_));
 AND3x1_ASAP7_75t_R _09173_ (.A(net4889),
    .B(_03145_),
    .C(net5063),
    .Y(_03152_));
 NOR2x1_ASAP7_75t_R _09174_ (.A(net5207),
    .B(_03149_),
    .Y(_03153_));
 NAND2x1_ASAP7_75t_R _09175_ (.A(net5064),
    .B(_03152_),
    .Y(_03154_));
 OA211x2_ASAP7_75t_R _09176_ (.A1(_03152_),
    .A2(_03153_),
    .B(_03154_),
    .C(net5362),
    .Y(_00740_));
 NOR2x1_ASAP7_75t_R _09177_ (.A(net5207),
    .B(_03151_),
    .Y(_03155_));
 INVx1_ASAP7_75t_R _09178_ (.A(_03155_),
    .Y(_03156_));
 OAI21x1_ASAP7_75t_R _09179_ (.A1(net5206),
    .A2(_03149_),
    .B(_03156_),
    .Y(_03157_));
 OA211x2_ASAP7_75t_R _09180_ (.A1(net5206),
    .A2(_03156_),
    .B(net5362),
    .C(_03157_),
    .Y(_00741_));
 INVx1_ASAP7_75t_R _09181_ (.A(_00538_),
    .Y(_03158_));
 AND5x1_ASAP7_75t_R _09182_ (.A(net4748),
    .B(_00110_),
    .C(net5153),
    .D(_03158_),
    .E(net4857),
    .Y(_03159_));
 AO21x1_ASAP7_75t_R _09183_ (.A1(_03159_),
    .A2(net4698),
    .B(net4699),
    .Y(_03160_));
 BUFx3_ASAP7_75t_R place2977 (.A(net2976),
    .Y(net2977));
 OA21x2_ASAP7_75t_R _09185_ (.A1(_03160_),
    .A2(net5199),
    .B(net5197),
    .Y(_03162_));
 NOR2x1_ASAP7_75t_R _09186_ (.A(net5360),
    .B(_03162_),
    .Y(_00743_));
 BUFx3_ASAP7_75t_R place2975 (.A(_06284_),
    .Y(net2975));
 NAND2x1_ASAP7_75t_R _09188_ (.A(net4974),
    .B(net5030),
    .Y(_03164_));
 INVx6_ASAP7_75t_R _09189_ (.A(net5198),
    .Y(_03165_));
 INVx1_ASAP7_75t_R _09190_ (.A(_00525_),
    .Y(_03166_));
 AND3x1_ASAP7_75t_R _09191_ (.A(_03166_),
    .B(net5176),
    .C(net5175),
    .Y(_03167_));
 INVx1_ASAP7_75t_R _09192_ (.A(_03167_),
    .Y(_03168_));
 NAND2x1_ASAP7_75t_R _09193_ (.A(net4680),
    .B(net4330),
    .Y(_03169_));
 XOR2x2_ASAP7_75t_R _09194_ (.A(_03169_),
    .B(net5174),
    .Y(_03170_));
 AO21x1_ASAP7_75t_R _09195_ (.A1(net4964),
    .A2(net5708),
    .B(net4971),
    .Y(_03171_));
 AND3x2_ASAP7_75t_R _09196_ (.A(_03171_),
    .B(net4973),
    .C(net4972),
    .Y(_03172_));
 XOR2x2_ASAP7_75t_R _09197_ (.A(_03172_),
    .B(net5196),
    .Y(_03173_));
 XOR2x2_ASAP7_75t_R _09198_ (.A(net4744),
    .B(net4973),
    .Y(_03174_));
 INVx1_ASAP7_75t_R _09199_ (.A(net4679),
    .Y(_03175_));
 XOR2x2_ASAP7_75t_R _09200_ (.A(net4841),
    .B(net4972),
    .Y(_03176_));
 INVx1_ASAP7_75t_R _09201_ (.A(net4732),
    .Y(_03177_));
 XOR2x2_ASAP7_75t_R _09202_ (.A(net4817),
    .B(net5173),
    .Y(_03178_));
 OR4x1_ASAP7_75t_R _09203_ (.A(net4967),
    .B(net4966),
    .C(_00531_),
    .D(_00527_),
    .Y(_03179_));
 INVx1_ASAP7_75t_R _09204_ (.A(_03179_),
    .Y(_03180_));
 AND5x1_ASAP7_75t_R _09205_ (.A(_03173_),
    .B(_03175_),
    .C(_03177_),
    .D(net4731),
    .E(_03180_),
    .Y(_03181_));
 OR3x1_ASAP7_75t_R _09206_ (.A(net4372),
    .B(net4373),
    .C(net4566),
    .Y(_03182_));
 XOR2x2_ASAP7_75t_R _09207_ (.A(net5195),
    .B(net4691),
    .Y(_03183_));
 INVx2_ASAP7_75t_R _09208_ (.A(_03183_),
    .Y(_03184_));
 XOR2x2_ASAP7_75t_R _09209_ (.A(_03182_),
    .B(net4565),
    .Y(_03185_));
 INVx1_ASAP7_75t_R _09210_ (.A(_03185_),
    .Y(_03186_));
 XOR2x2_ASAP7_75t_R _09211_ (.A(net4472),
    .B(net5182),
    .Y(_03187_));
 NAND2x1_ASAP7_75t_R _09212_ (.A(net4987),
    .B(net4986),
    .Y(_03188_));
 NOR2x1_ASAP7_75t_R _09213_ (.A(net5195),
    .B(net5196),
    .Y(_03189_));
 AND3x1_ASAP7_75t_R _09214_ (.A(_03189_),
    .B(net4977),
    .C(net4976),
    .Y(_03190_));
 AND5x1_ASAP7_75t_R _09215_ (.A(net4981),
    .B(_03190_),
    .C(net4980),
    .D(net4979),
    .E(net4978),
    .Y(_03191_));
 NOR2x1_ASAP7_75t_R _09216_ (.A(net5190),
    .B(net5191),
    .Y(_03192_));
 AND3x1_ASAP7_75t_R _09217_ (.A(_03192_),
    .B(net4985),
    .C(net4984),
    .Y(_03193_));
 AND3x1_ASAP7_75t_R _09218_ (.A(_03191_),
    .B(net4733),
    .C(_03193_),
    .Y(_03194_));
 INVx1_ASAP7_75t_R _09219_ (.A(_03194_),
    .Y(_03195_));
 NOR2x1_ASAP7_75t_R _09220_ (.A(_03188_),
    .B(_03195_),
    .Y(_03196_));
 INVx1_ASAP7_75t_R _09221_ (.A(_03196_),
    .Y(_03197_));
 OR5x1_ASAP7_75t_R _09222_ (.A(net5182),
    .B(_03197_),
    .C(net5183),
    .D(net5184),
    .E(net5185),
    .Y(_03198_));
 XOR2x2_ASAP7_75t_R _09223_ (.A(_03198_),
    .B(net4992),
    .Y(_03199_));
 INVx1_ASAP7_75t_R _09224_ (.A(_03199_),
    .Y(_03200_));
 NOR2x1_ASAP7_75t_R _09225_ (.A(_03187_),
    .B(_03200_),
    .Y(_03201_));
 OR3x1_ASAP7_75t_R _09226_ (.A(_02504_),
    .B(net5181),
    .C(net5182),
    .Y(_03202_));
 XOR2x2_ASAP7_75t_R _09227_ (.A(_03202_),
    .B(net5180),
    .Y(_03203_));
 INVx1_ASAP7_75t_R _09228_ (.A(_03203_),
    .Y(_03204_));
 AND2x2_ASAP7_75t_R _09229_ (.A(_03201_),
    .B(_03204_),
    .Y(_03205_));
 INVx1_ASAP7_75t_R _09230_ (.A(_03205_),
    .Y(_03206_));
 NOR2x1_ASAP7_75t_R _09231_ (.A(net5183),
    .B(net5184),
    .Y(_03207_));
 NOR2x1_ASAP7_75t_R _09232_ (.A(net5185),
    .B(net4524),
    .Y(_03208_));
 AOI21x1_ASAP7_75t_R _09233_ (.A1(net4989),
    .A2(_03208_),
    .B(net4990),
    .Y(_03209_));
 AOI21x1_ASAP7_75t_R _09234_ (.A1(_03207_),
    .A2(_03208_),
    .B(_03209_),
    .Y(_03210_));
 INVx1_ASAP7_75t_R _09235_ (.A(_03210_),
    .Y(_03211_));
 AND2x2_ASAP7_75t_R _09236_ (.A(net4729),
    .B(net4733),
    .Y(_03212_));
 XOR2x2_ASAP7_75t_R _09237_ (.A(_03212_),
    .B(net4982),
    .Y(_03213_));
 AND3x1_ASAP7_75t_R _09238_ (.A(_02497_),
    .B(net4978),
    .C(net4977),
    .Y(_03214_));
 AND2x2_ASAP7_75t_R _09239_ (.A(_03214_),
    .B(_02498_),
    .Y(_03215_));
 AND3x1_ASAP7_75t_R _09240_ (.A(_03215_),
    .B(net4982),
    .C(net4981),
    .Y(_03216_));
 XOR2x2_ASAP7_75t_R _09241_ (.A(_03216_),
    .B(net4983),
    .Y(_03217_));
 NOR2x1_ASAP7_75t_R _09242_ (.A(net4623),
    .B(_03217_),
    .Y(_03218_));
 INVx1_ASAP7_75t_R _09243_ (.A(_03218_),
    .Y(_03219_));
 AND2x4_ASAP7_75t_R _09244_ (.A(_03172_),
    .B(net4886),
    .Y(_03220_));
 AND3x2_ASAP7_75t_R _09245_ (.A(_03220_),
    .B(net4977),
    .C(net4976),
    .Y(_03221_));
 AND3x1_ASAP7_75t_R _09246_ (.A(_03221_),
    .B(net4979),
    .C(net4978),
    .Y(_03222_));
 XOR2x2_ASAP7_75t_R _09247_ (.A(_03222_),
    .B(net5193),
    .Y(_03223_));
 XOR2x2_ASAP7_75t_R _09248_ (.A(_03215_),
    .B(net5192),
    .Y(_03224_));
 AND2x4_ASAP7_75t_R _09249_ (.A(_03223_),
    .B(_03224_),
    .Y(_03225_));
 INVx2_ASAP7_75t_R _09250_ (.A(_03225_),
    .Y(_03226_));
 XOR2x2_ASAP7_75t_R _09251_ (.A(net4639),
    .B(net4977),
    .Y(_03227_));
 XOR2x2_ASAP7_75t_R _09252_ (.A(net4677),
    .B(net4976),
    .Y(_03228_));
 NOR2x1_ASAP7_75t_R _09253_ (.A(_03227_),
    .B(_03228_),
    .Y(_03229_));
 INVx1_ASAP7_75t_R _09254_ (.A(_03229_),
    .Y(_03230_));
 AND2x2_ASAP7_75t_R _09255_ (.A(net5176),
    .B(net5175),
    .Y(_03231_));
 AND4x1_ASAP7_75t_R _09256_ (.A(_03231_),
    .B(net5179),
    .C(net5709),
    .D(net5189),
    .Y(_03232_));
 AND3x1_ASAP7_75t_R _09257_ (.A(_03232_),
    .B(_00532_),
    .C(_03178_),
    .Y(_03233_));
 NOR2x1_ASAP7_75t_R _09258_ (.A(_03174_),
    .B(_03176_),
    .Y(_03234_));
 AND2x2_ASAP7_75t_R _09259_ (.A(_03233_),
    .B(_03234_),
    .Y(_03235_));
 INVx1_ASAP7_75t_R _09260_ (.A(_03173_),
    .Y(_03236_));
 NOR2x1_ASAP7_75t_R _09261_ (.A(_03184_),
    .B(_03236_),
    .Y(_03237_));
 AND2x2_ASAP7_75t_R _09262_ (.A(_03235_),
    .B(_03237_),
    .Y(_03238_));
 INVx2_ASAP7_75t_R _09263_ (.A(_03238_),
    .Y(_03239_));
 NOR2x1_ASAP7_75t_R _09264_ (.A(_03239_),
    .B(_03230_),
    .Y(_03240_));
 INVx1_ASAP7_75t_R _09265_ (.A(_03240_),
    .Y(_03241_));
 XOR2x2_ASAP7_75t_R _09266_ (.A(net4563),
    .B(net4979),
    .Y(_03242_));
 XOR2x2_ASAP7_75t_R _09267_ (.A(_03221_),
    .B(net4978),
    .Y(_03243_));
 NOR2x1_ASAP7_75t_R _09268_ (.A(_03242_),
    .B(_03243_),
    .Y(_03244_));
 INVx1_ASAP7_75t_R _09269_ (.A(_03244_),
    .Y(_03245_));
 OR3x2_ASAP7_75t_R _09270_ (.A(_03241_),
    .B(_03226_),
    .C(_03245_),
    .Y(_03246_));
 NOR2x1p5_ASAP7_75t_R _09271_ (.A(_03246_),
    .B(_03219_),
    .Y(_03247_));
 AND3x1_ASAP7_75t_R _09272_ (.A(net4729),
    .B(net4733),
    .C(net4885),
    .Y(_03248_));
 XOR2x2_ASAP7_75t_R _09273_ (.A(_03248_),
    .B(net4984),
    .Y(_03249_));
 INVx1_ASAP7_75t_R _09274_ (.A(_03249_),
    .Y(_03250_));
 OR3x1_ASAP7_75t_R _09275_ (.A(_02501_),
    .B(net5187),
    .C(net5188),
    .Y(_03251_));
 OR3x1_ASAP7_75t_R _09276_ (.A(_03251_),
    .B(net5185),
    .C(net5186),
    .Y(_03252_));
 XOR2x2_ASAP7_75t_R _09277_ (.A(_03252_),
    .B(net5184),
    .Y(_03253_));
 INVx1_ASAP7_75t_R _09278_ (.A(_03253_),
    .Y(_03254_));
 XOR2x2_ASAP7_75t_R _09279_ (.A(_03251_),
    .B(net5186),
    .Y(_03255_));
 XOR2x2_ASAP7_75t_R _09280_ (.A(net4564),
    .B(net4988),
    .Y(_03256_));
 NOR2x1_ASAP7_75t_R _09281_ (.A(_03255_),
    .B(_03256_),
    .Y(_03257_));
 AO21x1_ASAP7_75t_R _09282_ (.A1(_02500_),
    .A2(net4639),
    .B(net4985),
    .Y(_03258_));
 AND2x2_ASAP7_75t_R _09283_ (.A(_02502_),
    .B(_03258_),
    .Y(_03259_));
 XOR2x2_ASAP7_75t_R _09284_ (.A(net4678),
    .B(net4986),
    .Y(_03260_));
 NOR2x1_ASAP7_75t_R _09285_ (.A(_03259_),
    .B(_03260_),
    .Y(_03261_));
 AND2x2_ASAP7_75t_R _09286_ (.A(_03257_),
    .B(_03261_),
    .Y(_03262_));
 AND4x2_ASAP7_75t_R _09287_ (.A(_03247_),
    .B(_03250_),
    .C(_03254_),
    .D(_03262_),
    .Y(_03263_));
 NAND2x1p5_ASAP7_75t_R _09288_ (.A(_03263_),
    .B(_03211_),
    .Y(_03264_));
 OA21x2_ASAP7_75t_R _09289_ (.A1(_03264_),
    .A2(_03206_),
    .B(net4328),
    .Y(_03265_));
 OR3x1_ASAP7_75t_R _09290_ (.A(_03198_),
    .B(net5180),
    .C(net5181),
    .Y(_03266_));
 XOR2x2_ASAP7_75t_R _09291_ (.A(_03266_),
    .B(net5178),
    .Y(_03267_));
 XOR2x2_ASAP7_75t_R _09292_ (.A(net4365),
    .B(_03265_),
    .Y(_03268_));
 INVx1_ASAP7_75t_R _09293_ (.A(_03242_),
    .Y(_03269_));
 AND2x2_ASAP7_75t_R _09294_ (.A(net4522),
    .B(_03269_),
    .Y(_03270_));
 NOR2x1_ASAP7_75t_R _09295_ (.A(net4562),
    .B(_03243_),
    .Y(_03271_));
 INVx1_ASAP7_75t_R _09296_ (.A(_03228_),
    .Y(_03272_));
 NAND2x1_ASAP7_75t_R _09297_ (.A(_03183_),
    .B(_03272_),
    .Y(_03273_));
 INVx1_ASAP7_75t_R _09298_ (.A(net4731),
    .Y(_03274_));
 OR4x1_ASAP7_75t_R _09299_ (.A(net4732),
    .B(net4818),
    .C(_03274_),
    .D(_03168_),
    .Y(_03275_));
 OR4x1_ASAP7_75t_R _09300_ (.A(_03273_),
    .B(net4620),
    .C(net4679),
    .D(_03275_),
    .Y(_03276_));
 INVx1_ASAP7_75t_R _09301_ (.A(_03276_),
    .Y(_03277_));
 AND3x1_ASAP7_75t_R _09302_ (.A(_03270_),
    .B(net4519),
    .C(_03277_),
    .Y(_03278_));
 NOR2x1_ASAP7_75t_R _09303_ (.A(_03249_),
    .B(net4427),
    .Y(_03279_));
 INVx1_ASAP7_75t_R _09304_ (.A(_03213_),
    .Y(_03280_));
 AND2x2_ASAP7_75t_R _09305_ (.A(_03280_),
    .B(net4469),
    .Y(_03281_));
 AND3x1_ASAP7_75t_R _09306_ (.A(_03278_),
    .B(_03279_),
    .C(net4420),
    .Y(_03282_));
 NAND2x1_ASAP7_75t_R _09307_ (.A(net4366),
    .B(_03282_),
    .Y(_03283_));
 NOR2x1_ASAP7_75t_R _09308_ (.A(_03210_),
    .B(net4424),
    .Y(_03284_));
 NAND2x1_ASAP7_75t_R _09309_ (.A(_03284_),
    .B(net4325),
    .Y(_03285_));
 OAI21x1_ASAP7_75t_R _09310_ (.A1(_03283_),
    .A2(_03285_),
    .B(net4328),
    .Y(_03286_));
 XOR2x2_ASAP7_75t_R _09311_ (.A(_03286_),
    .B(net4369),
    .Y(_03287_));
 INVx1_ASAP7_75t_R _09312_ (.A(_03287_),
    .Y(_03288_));
 INVx1_ASAP7_75t_R _09313_ (.A(_02508_),
    .Y(_03289_));
 NOR2x1_ASAP7_75t_R _09314_ (.A(_03289_),
    .B(_03267_),
    .Y(_03290_));
 INVx1_ASAP7_75t_R _09315_ (.A(_03273_),
    .Y(_03291_));
 AND3x1_ASAP7_75t_R _09316_ (.A(_03271_),
    .B(_03181_),
    .C(_03291_),
    .Y(_03292_));
 AND3x1_ASAP7_75t_R _09317_ (.A(_03270_),
    .B(_03292_),
    .C(_03281_),
    .Y(_03293_));
 AND3x1_ASAP7_75t_R _09318_ (.A(_03293_),
    .B(_03279_),
    .C(net4422),
    .Y(_03294_));
 AND3x1_ASAP7_75t_R _09319_ (.A(_03294_),
    .B(net4423),
    .C(_03284_),
    .Y(_03295_));
 AND3x1_ASAP7_75t_R _09320_ (.A(_03290_),
    .B(_03205_),
    .C(_03295_),
    .Y(_03296_));
 NAND2x1_ASAP7_75t_R _09321_ (.A(_03265_),
    .B(_03296_),
    .Y(_03297_));
 AND3x1_ASAP7_75t_R _09322_ (.A(_03268_),
    .B(_03288_),
    .C(_03297_),
    .Y(_03298_));
 INVx2_ASAP7_75t_R _09323_ (.A(_03298_),
    .Y(_03299_));
 BUFx3_ASAP7_75t_R place2974 (.A(_06285_),
    .Y(net2974));
 NOR2x1_ASAP7_75t_R _09325_ (.A(_03289_),
    .B(_03263_),
    .Y(_03301_));
 XOR2x2_ASAP7_75t_R _09326_ (.A(_03301_),
    .B(net4324),
    .Y(_03302_));
 NOR2x1_ASAP7_75t_R _09327_ (.A(_03289_),
    .B(_03295_),
    .Y(_03303_));
 XNOR2x2_ASAP7_75t_R _09328_ (.A(net4428),
    .B(_03303_),
    .Y(_03304_));
 OAI21x1_ASAP7_75t_R _09329_ (.A1(net4428),
    .A2(net4084),
    .B(net4328),
    .Y(_03305_));
 XOR2x2_ASAP7_75t_R _09330_ (.A(_03305_),
    .B(net4370),
    .Y(_03306_));
 AND4x1_ASAP7_75t_R _09331_ (.A(_03297_),
    .B(_03302_),
    .C(_03304_),
    .D(_03306_),
    .Y(_03307_));
 AND3x1_ASAP7_75t_R _09332_ (.A(net4519),
    .B(net4566),
    .C(_03291_),
    .Y(_03308_));
 AND5x1_ASAP7_75t_R _09333_ (.A(_03279_),
    .B(_03308_),
    .C(net4420),
    .D(_03270_),
    .E(net4422),
    .Y(_03309_));
 AND5x1_ASAP7_75t_R _09334_ (.A(net4423),
    .B(_03290_),
    .C(_03284_),
    .D(_03205_),
    .E(_03309_),
    .Y(_03310_));
 NAND2x1_ASAP7_75t_R _09335_ (.A(net4040),
    .B(_03310_),
    .Y(_03311_));
 OAI21x1_ASAP7_75t_R _09336_ (.A1(_03299_),
    .A2(_03307_),
    .B(_03311_),
    .Y(_03312_));
 AND2x2_ASAP7_75t_R _09337_ (.A(_03283_),
    .B(net4328),
    .Y(_03313_));
 XOR2x2_ASAP7_75t_R _09338_ (.A(_03313_),
    .B(net4367),
    .Y(_03314_));
 INVx1_ASAP7_75t_R _09339_ (.A(net4520),
    .Y(_03315_));
 AND4x1_ASAP7_75t_R _09340_ (.A(net4468),
    .B(_03229_),
    .C(net4521),
    .D(net4621),
    .Y(_03316_));
 NOR2x1_ASAP7_75t_R _09341_ (.A(net4466),
    .B(_03249_),
    .Y(_03317_));
 NOR2x1_ASAP7_75t_R _09342_ (.A(net4619),
    .B(net4467),
    .Y(_03318_));
 AND5x1_ASAP7_75t_R _09343_ (.A(net4368),
    .B(_03316_),
    .C(net4426),
    .D(_03317_),
    .E(_03318_),
    .Y(_03319_));
 AND3x1_ASAP7_75t_R _09344_ (.A(_03319_),
    .B(net4676),
    .C(_03315_),
    .Y(_03320_));
 AOI21x1_ASAP7_75t_R _09345_ (.A1(net4676),
    .A2(_03319_),
    .B(_03315_),
    .Y(_03321_));
 OA21x2_ASAP7_75t_R _09346_ (.A1(_03320_),
    .A2(_03321_),
    .B(net4329),
    .Y(_03322_));
 AO21x1_ASAP7_75t_R _09347_ (.A1(net4275),
    .A2(_03315_),
    .B(_03322_),
    .Y(_03323_));
 NAND2x1_ASAP7_75t_R _09348_ (.A(_03314_),
    .B(_03323_),
    .Y(_03324_));
 INVx1_ASAP7_75t_R _09349_ (.A(net4040),
    .Y(_03325_));
 INVx1_ASAP7_75t_R _09350_ (.A(_03304_),
    .Y(_03326_));
 AO21x2_ASAP7_75t_R _09351_ (.A1(_03296_),
    .A2(_03265_),
    .B(_03326_),
    .Y(_03327_));
 INVx1_ASAP7_75t_R _09352_ (.A(_03327_),
    .Y(_03328_));
 NAND2x1_ASAP7_75t_R _09353_ (.A(_03325_),
    .B(_03328_),
    .Y(_03329_));
 AOI21x1_ASAP7_75t_R _09354_ (.A1(_03325_),
    .A2(_03324_),
    .B(_03327_),
    .Y(_03330_));
 OAI21x1_ASAP7_75t_R _09355_ (.A1(net4083),
    .A2(_03329_),
    .B(_03330_),
    .Y(_03331_));
 INVx1_ASAP7_75t_R _09356_ (.A(_03306_),
    .Y(_03332_));
 NAND2x1_ASAP7_75t_R _09357_ (.A(_03332_),
    .B(net4014),
    .Y(_03333_));
 INVx1_ASAP7_75t_R _09358_ (.A(_03333_),
    .Y(_03334_));
 XOR2x2_ASAP7_75t_R _09359_ (.A(_03331_),
    .B(_03334_),
    .Y(_03335_));
 NOR2x1_ASAP7_75t_R _09360_ (.A(net3982),
    .B(net3983),
    .Y(_03336_));
 AOI21x1_ASAP7_75t_R _09361_ (.A1(net3983),
    .A2(_03335_),
    .B(_03336_),
    .Y(_03337_));
 NOR2x1_ASAP7_75t_R _09362_ (.A(net3989),
    .B(net3997),
    .Y(_03338_));
 NOR2x1_ASAP7_75t_R _09363_ (.A(net4150),
    .B(_03338_),
    .Y(_03339_));
 AND2x4_ASAP7_75t_R _09364_ (.A(_03337_),
    .B(_03339_),
    .Y(_03340_));
 INVx1_ASAP7_75t_R _09365_ (.A(_03338_),
    .Y(_03341_));
 AND2x2_ASAP7_75t_R _09366_ (.A(_03268_),
    .B(net4014),
    .Y(_03342_));
 AND2x2_ASAP7_75t_R _09367_ (.A(_03341_),
    .B(_03342_),
    .Y(_03343_));
 NOR2x1_ASAP7_75t_R _09368_ (.A(_03312_),
    .B(net4013),
    .Y(_03344_));
 INVx1_ASAP7_75t_R _09369_ (.A(_03312_),
    .Y(_03345_));
 NOR2x1_ASAP7_75t_R _09370_ (.A(net4041),
    .B(_03345_),
    .Y(_03346_));
 OAI21x1_ASAP7_75t_R _09371_ (.A1(_03346_),
    .A2(_03344_),
    .B(net4149),
    .Y(_03347_));
 NOR2x2_ASAP7_75t_R _09372_ (.A(_03347_),
    .B(net4012),
    .Y(_03348_));
 INVx2_ASAP7_75t_R _09373_ (.A(_03348_),
    .Y(_03349_));
 OA21x2_ASAP7_75t_R _09374_ (.A1(_03340_),
    .A2(_03343_),
    .B(_03349_),
    .Y(_03350_));
 XNOR2x2_ASAP7_75t_R _09375_ (.A(net3962),
    .B(_03350_),
    .Y(_03351_));
 NAND2x1_ASAP7_75t_R _09376_ (.A(net4041),
    .B(net3984),
    .Y(_03352_));
 XOR2x2_ASAP7_75t_R _09377_ (.A(_03352_),
    .B(net3996),
    .Y(_03353_));
 AOI21x1_ASAP7_75t_R _09378_ (.A1(_03340_),
    .A2(_03349_),
    .B(_03343_),
    .Y(_03354_));
 INVx2_ASAP7_75t_R _09379_ (.A(_03354_),
    .Y(_03355_));
 XOR2x2_ASAP7_75t_R _09380_ (.A(_03353_),
    .B(net3951),
    .Y(_03356_));
 NAND2x1_ASAP7_75t_R _09381_ (.A(_03356_),
    .B(_03355_),
    .Y(_03357_));
 OAI21x1_ASAP7_75t_R _09382_ (.A1(net3961),
    .A2(_03355_),
    .B(_03357_),
    .Y(_03358_));
 NOR2x2_ASAP7_75t_R _09383_ (.A(_03358_),
    .B(_03351_),
    .Y(_03359_));
 AND2x2_ASAP7_75t_R _09384_ (.A(_03350_),
    .B(net3962),
    .Y(_03360_));
 INVx1_ASAP7_75t_R _09385_ (.A(_03340_),
    .Y(_03361_));
 NOR2x1_ASAP7_75t_R _09386_ (.A(net3945),
    .B(_03361_),
    .Y(_03362_));
 INVx1_ASAP7_75t_R _09387_ (.A(_03362_),
    .Y(_03363_));
 OA21x2_ASAP7_75t_R _09388_ (.A1(_03360_),
    .A2(net3970),
    .B(_03363_),
    .Y(_03364_));
 INVx1_ASAP7_75t_R _09389_ (.A(_03344_),
    .Y(_03365_));
 INVx1_ASAP7_75t_R _09390_ (.A(_03346_),
    .Y(_03366_));
 NAND2x1_ASAP7_75t_R _09391_ (.A(_03365_),
    .B(_03366_),
    .Y(_03367_));
 NAND2x1p5_ASAP7_75t_R _09392_ (.A(net4149),
    .B(net5673),
    .Y(_03368_));
 NOR2x1p5_ASAP7_75t_R _09393_ (.A(net4149),
    .B(_03354_),
    .Y(_03369_));
 INVx2_ASAP7_75t_R _09394_ (.A(_03369_),
    .Y(_03370_));
 INVx1_ASAP7_75t_R _09395_ (.A(net4148),
    .Y(_03371_));
 AOI21x1_ASAP7_75t_R _09396_ (.A1(_03370_),
    .A2(_03368_),
    .B(_03371_),
    .Y(_03372_));
 NAND2x2_ASAP7_75t_R _09397_ (.A(_03372_),
    .B(net3944),
    .Y(_03373_));
 OAI21x1_ASAP7_75t_R _09398_ (.A1(_03359_),
    .A2(_03364_),
    .B(_03373_),
    .Y(_03374_));
 XOR2x2_ASAP7_75t_R _09399_ (.A(_03374_),
    .B(net3890),
    .Y(_03375_));
 NAND2x1_ASAP7_75t_R _09400_ (.A(net3878),
    .B(net3876),
    .Y(_03376_));
 OAI21x1_ASAP7_75t_R _09401_ (.A1(net3890),
    .A2(net3870),
    .B(net3914),
    .Y(_03377_));
 NAND2x2_ASAP7_75t_R _09402_ (.A(_03377_),
    .B(_03376_),
    .Y(_03378_));
 INVx1_ASAP7_75t_R _09403_ (.A(_03375_),
    .Y(_03379_));
 NAND2x1_ASAP7_75t_R _09404_ (.A(net3913),
    .B(net3903),
    .Y(_03380_));
 INVx1_ASAP7_75t_R _09405_ (.A(_03380_),
    .Y(_03381_));
 INVx1_ASAP7_75t_R _09406_ (.A(net3912),
    .Y(_03382_));
 OAI21x1_ASAP7_75t_R _09407_ (.A1(net3911),
    .A2(_03382_),
    .B(net3944),
    .Y(_03383_));
 AOI211x1_ASAP7_75t_R _09408_ (.A1(net3877),
    .A2(_03383_),
    .B(net3904),
    .C(net4082),
    .Y(_03384_));
 AOI21x1_ASAP7_75t_R _09409_ (.A1(_03359_),
    .A2(_03373_),
    .B(_03364_),
    .Y(_03385_));
 NOR2x1_ASAP7_75t_R _09410_ (.A(_03385_),
    .B(net4148),
    .Y(_03386_));
 NOR2x1_ASAP7_75t_R _09411_ (.A(net4276),
    .B(_03294_),
    .Y(_03387_));
 XNOR2x2_ASAP7_75t_R _09412_ (.A(net4467),
    .B(_03387_),
    .Y(_03388_));
 OAI21x1_ASAP7_75t_R _09413_ (.A1(_03384_),
    .A2(_03386_),
    .B(net4146),
    .Y(_03389_));
 NOR2x1p5_ASAP7_75t_R _09414_ (.A(_03389_),
    .B(_03381_),
    .Y(_03390_));
 NOR2x1_ASAP7_75t_R _09415_ (.A(net3951),
    .B(net3921),
    .Y(_03391_));
 INVx1_ASAP7_75t_R _09416_ (.A(net4149),
    .Y(_03392_));
 INVx1_ASAP7_75t_R _09417_ (.A(_03367_),
    .Y(_03393_));
 OA21x2_ASAP7_75t_R _09418_ (.A1(net3921),
    .A2(_03392_),
    .B(_03393_),
    .Y(_03394_));
 NOR2x1_ASAP7_75t_R _09419_ (.A(_03391_),
    .B(_03394_),
    .Y(_03395_));
 XNOR2x2_ASAP7_75t_R _09420_ (.A(net3889),
    .B(_03395_),
    .Y(_03396_));
 NAND2x2_ASAP7_75t_R _09421_ (.A(net3902),
    .B(net5695),
    .Y(_03397_));
 OAI21x1_ASAP7_75t_R _09422_ (.A1(net5683),
    .A2(_03396_),
    .B(_03397_),
    .Y(_03398_));
 AOI211x1_ASAP7_75t_R _09423_ (.A1(net5697),
    .A2(_03379_),
    .B(_03390_),
    .C(net3845),
    .Y(_03399_));
 NOR2x2_ASAP7_75t_R _09424_ (.A(_03379_),
    .B(_03398_),
    .Y(_03400_));
 NAND2x1p5_ASAP7_75t_R _09425_ (.A(net4148),
    .B(net5696),
    .Y(_03401_));
 NOR2x1_ASAP7_75t_R _09426_ (.A(net4082),
    .B(_03383_),
    .Y(_03402_));
 INVx1_ASAP7_75t_R _09427_ (.A(_03359_),
    .Y(_03403_));
 INVx1_ASAP7_75t_R _09428_ (.A(_03364_),
    .Y(_03404_));
 OAI21x1_ASAP7_75t_R _09429_ (.A1(_03402_),
    .A2(_03403_),
    .B(_03404_),
    .Y(_03405_));
 NAND2x1_ASAP7_75t_R _09430_ (.A(_03405_),
    .B(net4082),
    .Y(_03406_));
 INVx1_ASAP7_75t_R _09431_ (.A(_03388_),
    .Y(_03407_));
 AOI21x1_ASAP7_75t_R _09432_ (.A1(_03401_),
    .A2(_03406_),
    .B(_03407_),
    .Y(_03408_));
 NAND2x1p5_ASAP7_75t_R _09433_ (.A(net3888),
    .B(_03408_),
    .Y(_03409_));
 NAND2x2_ASAP7_75t_R _09434_ (.A(net3828),
    .B(net3817),
    .Y(_03410_));
 OAI21x1_ASAP7_75t_R _09435_ (.A1(net3859),
    .A2(_03399_),
    .B(_03410_),
    .Y(_03411_));
 NAND2x1_ASAP7_75t_R _09436_ (.A(net3858),
    .B(net3844),
    .Y(_03412_));
 INVx1_ASAP7_75t_R _09437_ (.A(net3825),
    .Y(_03413_));
 NOR2x1_ASAP7_75t_R _09438_ (.A(net3876),
    .B(net3887),
    .Y(_03414_));
 AOI21x1_ASAP7_75t_R _09439_ (.A1(net3889),
    .A2(net3857),
    .B(net3902),
    .Y(_03415_));
 OAI21x1_ASAP7_75t_R _09440_ (.A1(_03414_),
    .A2(_03415_),
    .B(net3859),
    .Y(_03416_));
 OAI21x1_ASAP7_75t_R _09441_ (.A1(_03416_),
    .A2(_03390_),
    .B(net3847),
    .Y(_03417_));
 NOR2x1_ASAP7_75t_R _09442_ (.A(net4081),
    .B(_03417_),
    .Y(_03418_));
 INVx1_ASAP7_75t_R _09443_ (.A(net5697),
    .Y(_03419_));
 AOI21x1_ASAP7_75t_R _09444_ (.A1(_03409_),
    .A2(_03400_),
    .B(_03419_),
    .Y(_03420_));
 NOR2x1_ASAP7_75t_R _09445_ (.A(net4147),
    .B(_03420_),
    .Y(_03421_));
 AOI21x1_ASAP7_75t_R _09446_ (.A1(net4418),
    .A2(net4219),
    .B(net4276),
    .Y(_03422_));
 XNOR2x2_ASAP7_75t_R _09447_ (.A(net4619),
    .B(_03422_),
    .Y(_03423_));
 OAI21x1_ASAP7_75t_R _09448_ (.A1(_03418_),
    .A2(_03421_),
    .B(net4080),
    .Y(_03424_));
 NOR2x1_ASAP7_75t_R _09449_ (.A(net3816),
    .B(_03424_),
    .Y(_03425_));
 NOR2x1_ASAP7_75t_R _09450_ (.A(net3848),
    .B(net3817),
    .Y(_03426_));
 XOR2x2_ASAP7_75t_R _09451_ (.A(_03380_),
    .B(net4082),
    .Y(_03427_));
 NAND2x2_ASAP7_75t_R _09452_ (.A(net3888),
    .B(net3869),
    .Y(_03428_));
 OAI21x1_ASAP7_75t_R _09453_ (.A1(net3869),
    .A2(_03427_),
    .B(_03428_),
    .Y(_03429_));
 AOI21x1_ASAP7_75t_R _09454_ (.A1(net3827),
    .A2(_03417_),
    .B(_03429_),
    .Y(_03430_));
 NOR2x1_ASAP7_75t_R _09455_ (.A(_03426_),
    .B(_03430_),
    .Y(_03431_));
 OAI21x1_ASAP7_75t_R _09456_ (.A1(net3791),
    .A2(_03425_),
    .B(net3790),
    .Y(_03432_));
 INVx8_ASAP7_75t_R _09457_ (.A(net6002),
    .Y(_03433_));
 OA21x2_ASAP7_75t_R _09458_ (.A1(_03390_),
    .A2(net5697),
    .B(net3845),
    .Y(_03434_));
 NOR2x2_ASAP7_75t_R _09459_ (.A(_03399_),
    .B(_03434_),
    .Y(_03435_));
 INVx2_ASAP7_75t_R _09460_ (.A(net6001),
    .Y(_03436_));
 NOR2x2_ASAP7_75t_R _09461_ (.A(_03436_),
    .B(_03433_),
    .Y(_03437_));
 NAND2x1_ASAP7_75t_R _09462_ (.A(_03417_),
    .B(net4081),
    .Y(_03438_));
 NAND2x1p5_ASAP7_75t_R _09463_ (.A(_03420_),
    .B(net4147),
    .Y(_03439_));
 INVx1_ASAP7_75t_R _09464_ (.A(_03423_),
    .Y(_03440_));
 AOI21x1_ASAP7_75t_R _09465_ (.A1(_03438_),
    .A2(_03439_),
    .B(_03440_),
    .Y(_03441_));
 AOI21x1_ASAP7_75t_R _09466_ (.A1(net3826),
    .A2(_03441_),
    .B(_03431_),
    .Y(_03442_));
 OAI21x1_ASAP7_75t_R _09467_ (.A1(_03433_),
    .A2(_03437_),
    .B(_03442_),
    .Y(_03443_));
 NAND2x1_ASAP7_75t_R _09468_ (.A(_03432_),
    .B(_03443_),
    .Y(_03444_));
 OAI21x1_ASAP7_75t_R _09469_ (.A1(_03430_),
    .A2(_03426_),
    .B(_03435_),
    .Y(_03445_));
 AOI21x1_ASAP7_75t_R _09470_ (.A1(net3826),
    .A2(_03441_),
    .B(_03445_),
    .Y(_03446_));
 AO21x2_ASAP7_75t_R _09471_ (.A1(net3753),
    .A2(net3789),
    .B(_03446_),
    .Y(_03447_));
 OAI21x1_ASAP7_75t_R _09472_ (.A1(_03425_),
    .A2(net3787),
    .B(net3791),
    .Y(_03448_));
 NOR2x1_ASAP7_75t_R _09473_ (.A(_03413_),
    .B(_03417_),
    .Y(_03449_));
 XOR2x2_ASAP7_75t_R _09474_ (.A(_03412_),
    .B(net4081),
    .Y(_03450_));
 NOR2x1_ASAP7_75t_R _09475_ (.A(_03450_),
    .B(_03420_),
    .Y(_03451_));
 NOR2x2_ASAP7_75t_R _09476_ (.A(_03449_),
    .B(_03451_),
    .Y(_03452_));
 INVx2_ASAP7_75t_R _09477_ (.A(_03452_),
    .Y(_03453_));
 AOI21x1_ASAP7_75t_R _09478_ (.A1(net3768),
    .A2(_03448_),
    .B(net3759),
    .Y(_03454_));
 NOR2x1_ASAP7_75t_R _09479_ (.A(_03453_),
    .B(_03445_),
    .Y(_03455_));
 OAI21x1_ASAP7_75t_R _09480_ (.A1(net3769),
    .A2(_03455_),
    .B(net3768),
    .Y(_03456_));
 NOR2x1_ASAP7_75t_R _09481_ (.A(net3767),
    .B(_03456_),
    .Y(_03457_));
 NOR2x1_ASAP7_75t_R _09482_ (.A(_03454_),
    .B(_03457_),
    .Y(_03458_));
 INVx2_ASAP7_75t_R _09483_ (.A(_03458_),
    .Y(_03459_));
 NOR2x1_ASAP7_75t_R _09484_ (.A(net4276),
    .B(_03282_),
    .Y(_03460_));
 INVx1_ASAP7_75t_R _09485_ (.A(net4466),
    .Y(_03461_));
 XOR2x2_ASAP7_75t_R _09486_ (.A(_03460_),
    .B(_03461_),
    .Y(_03462_));
 OAI21x1_ASAP7_75t_R _09487_ (.A1(net3770),
    .A2(_03446_),
    .B(net4039),
    .Y(_03463_));
 INVx1_ASAP7_75t_R _09488_ (.A(_03445_),
    .Y(_03464_));
 NAND2x1_ASAP7_75t_R _09489_ (.A(net3826),
    .B(_03441_),
    .Y(_03465_));
 AOI21x1_ASAP7_75t_R _09490_ (.A1(_03465_),
    .A2(_03464_),
    .B(_03433_),
    .Y(_03466_));
 NAND2x2_ASAP7_75t_R _09491_ (.A(net4080),
    .B(_03466_),
    .Y(_03467_));
 NAND2x1_ASAP7_75t_R _09492_ (.A(net3803),
    .B(net3788),
    .Y(_03468_));
 INVx1_ASAP7_75t_R _09493_ (.A(_03468_),
    .Y(_03469_));
 AOI21x1_ASAP7_75t_R _09494_ (.A1(_03463_),
    .A2(_03467_),
    .B(_03469_),
    .Y(_03470_));
 NAND2x1p5_ASAP7_75t_R _09495_ (.A(_03470_),
    .B(_03462_),
    .Y(_03471_));
 NAND2x1_ASAP7_75t_R _09496_ (.A(_03459_),
    .B(net3713),
    .Y(_03472_));
 AO21x1_ASAP7_75t_R _09497_ (.A1(net3739),
    .A2(net3740),
    .B(_03472_),
    .Y(_03473_));
 INVx1_ASAP7_75t_R _09498_ (.A(_03462_),
    .Y(_03474_));
 INVx2_ASAP7_75t_R _09499_ (.A(_03470_),
    .Y(_03475_));
 NAND2x1_ASAP7_75t_R _09500_ (.A(net3767),
    .B(_03456_),
    .Y(_03476_));
 INVx1_ASAP7_75t_R _09501_ (.A(_03429_),
    .Y(_03477_));
 NOR2x1_ASAP7_75t_R _09502_ (.A(_03477_),
    .B(net3815),
    .Y(_03478_));
 XOR2x2_ASAP7_75t_R _09503_ (.A(_03429_),
    .B(net3846),
    .Y(_03479_));
 NOR2x1_ASAP7_75t_R _09504_ (.A(_03479_),
    .B(net3804),
    .Y(_03480_));
 NOR2x1_ASAP7_75t_R _09505_ (.A(_03478_),
    .B(_03480_),
    .Y(_03481_));
 NAND3x1_ASAP7_75t_R _09506_ (.A(_03481_),
    .B(_03452_),
    .C(net6001),
    .Y(_03482_));
 AOI21x1_ASAP7_75t_R _09507_ (.A1(_03482_),
    .A2(net3791),
    .B(net3771),
    .Y(_03483_));
 NAND2x1_ASAP7_75t_R _09508_ (.A(net3759),
    .B(_03483_),
    .Y(_03484_));
 AOI21x1_ASAP7_75t_R _09509_ (.A1(_03476_),
    .A2(_03484_),
    .B(_03444_),
    .Y(_03485_));
 OAI21x1_ASAP7_75t_R _09510_ (.A1(_03474_),
    .A2(_03475_),
    .B(_03485_),
    .Y(_03486_));
 INVx1_ASAP7_75t_R _09511_ (.A(net3702),
    .Y(_03487_));
 AOI21x1_ASAP7_75t_R _09512_ (.A1(_03473_),
    .A2(net3740),
    .B(_03487_),
    .Y(_03488_));
 INVx3_ASAP7_75t_R _09513_ (.A(_03447_),
    .Y(_03489_));
 AOI211x1_ASAP7_75t_R _09514_ (.A1(_03485_),
    .A2(_03475_),
    .B(_03489_),
    .C(_03474_),
    .Y(_03490_));
 AOI21x1_ASAP7_75t_R _09515_ (.A1(net3739),
    .A2(_03486_),
    .B(net4145),
    .Y(_03491_));
 NAND2x1_ASAP7_75t_R _09516_ (.A(_03463_),
    .B(_03467_),
    .Y(_03492_));
 OAI21x1_ASAP7_75t_R _09517_ (.A1(_03491_),
    .A2(_03490_),
    .B(net3719),
    .Y(_03493_));
 INVx1_ASAP7_75t_R _09518_ (.A(_03493_),
    .Y(_03494_));
 NOR2x1_ASAP7_75t_R _09519_ (.A(net4276),
    .B(net4219),
    .Y(_03495_));
 XOR2x2_ASAP7_75t_R _09520_ (.A(_03495_),
    .B(net4560),
    .Y(_03496_));
 NAND2x1_ASAP7_75t_R _09521_ (.A(net4080),
    .B(_03448_),
    .Y(_03497_));
 AOI21x1_ASAP7_75t_R _09522_ (.A1(_03469_),
    .A2(_03497_),
    .B(net3752),
    .Y(_03498_));
 AND4x1_ASAP7_75t_R _09523_ (.A(_03489_),
    .B(_03498_),
    .C(net4145),
    .D(_03492_),
    .Y(_03499_));
 INVx1_ASAP7_75t_R _09524_ (.A(_03492_),
    .Y(_03500_));
 NOR2x1_ASAP7_75t_R _09525_ (.A(_03474_),
    .B(_03500_),
    .Y(_03501_));
 INVx2_ASAP7_75t_R _09526_ (.A(net5706),
    .Y(_03502_));
 OAI21x1_ASAP7_75t_R _09527_ (.A1(_03454_),
    .A2(_03457_),
    .B(_03502_),
    .Y(_03503_));
 OAI21x1_ASAP7_75t_R _09528_ (.A1(_03498_),
    .A2(_03503_),
    .B(net3739),
    .Y(_03504_));
 AOI21x1_ASAP7_75t_R _09529_ (.A1(_03501_),
    .A2(_03504_),
    .B(net5699),
    .Y(_03505_));
 NOR2x1p5_ASAP7_75t_R _09530_ (.A(_03499_),
    .B(_03505_),
    .Y(_03506_));
 AO21x1_ASAP7_75t_R _09531_ (.A1(_03494_),
    .A2(_03496_),
    .B(_03506_),
    .Y(_03507_));
 OAI21x1_ASAP7_75t_R _09532_ (.A1(_03489_),
    .A2(_03485_),
    .B(_03471_),
    .Y(_03508_));
 XOR2x2_ASAP7_75t_R _09533_ (.A(_03459_),
    .B(_03508_),
    .Y(_03509_));
 NAND2x1_ASAP7_75t_R _09534_ (.A(net3690),
    .B(_03507_),
    .Y(_03510_));
 OAI21x1_ASAP7_75t_R _09535_ (.A1(net3661),
    .A2(_03507_),
    .B(_03510_),
    .Y(_03511_));
 INVx2_ASAP7_75t_R _09536_ (.A(_03488_),
    .Y(_03512_));
 INVx2_ASAP7_75t_R _09537_ (.A(_03509_),
    .Y(_03513_));
 INVx2_ASAP7_75t_R _09538_ (.A(_03506_),
    .Y(_03514_));
 NAND2x1p5_ASAP7_75t_R _09539_ (.A(_03514_),
    .B(_03513_),
    .Y(_03515_));
 INVx1_ASAP7_75t_R _09540_ (.A(_03496_),
    .Y(_03516_));
 NOR2x1p5_ASAP7_75t_R _09541_ (.A(_03493_),
    .B(_03516_),
    .Y(_03517_));
 AOI21x1_ASAP7_75t_R _09542_ (.A1(_03512_),
    .A2(_03515_),
    .B(_03517_),
    .Y(_03518_));
 XOR2x2_ASAP7_75t_R _09543_ (.A(net3660),
    .B(_03518_),
    .Y(_03519_));
 NOR2x2_ASAP7_75t_R _09544_ (.A(_03509_),
    .B(_03506_),
    .Y(_03520_));
 OAI21x1_ASAP7_75t_R _09545_ (.A1(net3701),
    .A2(_03491_),
    .B(_03496_),
    .Y(_03521_));
 NOR2x2_ASAP7_75t_R _09546_ (.A(net3721),
    .B(net3710),
    .Y(_03522_));
 OAI21x1_ASAP7_75t_R _09547_ (.A1(net3720),
    .A2(_03522_),
    .B(net4145),
    .Y(_03523_));
 INVx1_ASAP7_75t_R _09548_ (.A(_03501_),
    .Y(_03524_));
 INVx1_ASAP7_75t_R _09549_ (.A(net5699),
    .Y(_03525_));
 AOI21x1_ASAP7_75t_R _09550_ (.A1(_03525_),
    .A2(net3712),
    .B(net3720),
    .Y(_03526_));
 NOR2x1_ASAP7_75t_R _09551_ (.A(_03524_),
    .B(_03526_),
    .Y(_03527_));
 AOI21x1_ASAP7_75t_R _09552_ (.A1(net3711),
    .A2(_03523_),
    .B(_03527_),
    .Y(_03528_));
 INVx1_ASAP7_75t_R _09553_ (.A(_03528_),
    .Y(_03529_));
 AOI211x1_ASAP7_75t_R _09554_ (.A1(_03520_),
    .A2(net3672),
    .B(_03529_),
    .C(net3661),
    .Y(_03530_));
 OAI21x1_ASAP7_75t_R _09555_ (.A1(net4038),
    .A2(net5698),
    .B(_03520_),
    .Y(_03531_));
 XOR2x2_ASAP7_75t_R _09556_ (.A(_03521_),
    .B(_03528_),
    .Y(_03532_));
 AOI21x1_ASAP7_75t_R _09557_ (.A1(_03512_),
    .A2(_03531_),
    .B(_03532_),
    .Y(_03533_));
 NOR2x1_ASAP7_75t_R _09558_ (.A(_03530_),
    .B(_03533_),
    .Y(_03534_));
 NAND2x2_ASAP7_75t_R _09559_ (.A(_03534_),
    .B(_03519_),
    .Y(_03535_));
 INVx1_ASAP7_75t_R _09560_ (.A(net3701),
    .Y(_03536_));
 INVx1_ASAP7_75t_R _09561_ (.A(_03491_),
    .Y(_03537_));
 NAND2x1_ASAP7_75t_R _09562_ (.A(_03536_),
    .B(_03537_),
    .Y(_03538_));
 INVx1_ASAP7_75t_R _09563_ (.A(net3658),
    .Y(_03539_));
 OA21x2_ASAP7_75t_R _09564_ (.A1(_03520_),
    .A2(net3661),
    .B(net4038),
    .Y(_03540_));
 AOI211x1_ASAP7_75t_R _09565_ (.A1(_03520_),
    .A2(_03493_),
    .B(net4038),
    .C(net3661),
    .Y(_03541_));
 OR3x1_ASAP7_75t_R _09566_ (.A(_03293_),
    .B(net4373),
    .C(net4372),
    .Y(_03542_));
 XOR2x2_ASAP7_75t_R _09567_ (.A(_03542_),
    .B(net4427),
    .Y(_03543_));
 OAI21x1_ASAP7_75t_R _09568_ (.A1(_03541_),
    .A2(_03540_),
    .B(_03543_),
    .Y(_03544_));
 NOR2x1p5_ASAP7_75t_R _09569_ (.A(_03539_),
    .B(_03544_),
    .Y(_03545_));
 AOI21x1_ASAP7_75t_R _09570_ (.A1(net3612),
    .A2(net3600),
    .B(net3607),
    .Y(_03546_));
 INVx1_ASAP7_75t_R _09571_ (.A(net3608),
    .Y(_03547_));
 XOR2x2_ASAP7_75t_R _09572_ (.A(_03546_),
    .B(_03547_),
    .Y(_03548_));
 OAI21x1_ASAP7_75t_R _09573_ (.A1(_03517_),
    .A2(_03515_),
    .B(net3650),
    .Y(_03549_));
 XOR2x2_ASAP7_75t_R _09574_ (.A(_03538_),
    .B(net4079),
    .Y(_03550_));
 NAND2x1_ASAP7_75t_R _09575_ (.A(_03550_),
    .B(_03549_),
    .Y(_03551_));
 OAI21x1_ASAP7_75t_R _09576_ (.A1(_03539_),
    .A2(net3634),
    .B(_03551_),
    .Y(_03552_));
 INVx1_ASAP7_75t_R _09577_ (.A(net3599),
    .Y(_03553_));
 OAI21x1_ASAP7_75t_R _09578_ (.A1(_03535_),
    .A2(_03545_),
    .B(_03511_),
    .Y(_03554_));
 XNOR2x2_ASAP7_75t_R _09579_ (.A(_03552_),
    .B(net3635),
    .Y(_03555_));
 NAND2x1_ASAP7_75t_R _09580_ (.A(_03555_),
    .B(_03554_),
    .Y(_03556_));
 OAI21x1_ASAP7_75t_R _09581_ (.A1(_03553_),
    .A2(net3593),
    .B(_03556_),
    .Y(_03557_));
 NOR2x2_ASAP7_75t_R _09582_ (.A(_03548_),
    .B(_03557_),
    .Y(_03558_));
 NOR2x1_ASAP7_75t_R _09583_ (.A(net3649),
    .B(net5689),
    .Y(_03559_));
 INVx1_ASAP7_75t_R _09584_ (.A(net3632),
    .Y(_03560_));
 INVx1_ASAP7_75t_R _09585_ (.A(net4274),
    .Y(_03561_));
 NAND2x2_ASAP7_75t_R _09586_ (.A(_03561_),
    .B(_03554_),
    .Y(_03562_));
 OAI21x1_ASAP7_75t_R _09587_ (.A1(net5689),
    .A2(net3649),
    .B(net3659),
    .Y(_03563_));
 NAND3x1_ASAP7_75t_R _09588_ (.A(net3610),
    .B(net3608),
    .C(_03563_),
    .Y(_03564_));
 NAND3x1_ASAP7_75t_R _09589_ (.A(_03564_),
    .B(net4274),
    .C(_03511_),
    .Y(_03565_));
 NAND2x1_ASAP7_75t_R _09590_ (.A(net4277),
    .B(net4330),
    .Y(_03566_));
 XOR2x2_ASAP7_75t_R _09591_ (.A(_03566_),
    .B(net4623),
    .Y(_03567_));
 INVx1_ASAP7_75t_R _09592_ (.A(_03567_),
    .Y(_03568_));
 AOI21x1_ASAP7_75t_R _09593_ (.A1(_03562_),
    .A2(_03565_),
    .B(_03568_),
    .Y(_03569_));
 NAND2x1p5_ASAP7_75t_R _09594_ (.A(_03569_),
    .B(_03560_),
    .Y(_03570_));
 NOR2x1_ASAP7_75t_R _09595_ (.A(_03547_),
    .B(net3607),
    .Y(_03571_));
 NAND2x1_ASAP7_75t_R _09596_ (.A(net3611),
    .B(_03571_),
    .Y(_03572_));
 AO21x1_ASAP7_75t_R _09597_ (.A1(_03554_),
    .A2(_03571_),
    .B(net3611),
    .Y(_03573_));
 NAND2x1p5_ASAP7_75t_R _09598_ (.A(_03573_),
    .B(_03572_),
    .Y(_03574_));
 INVx4_ASAP7_75t_R _09599_ (.A(_03574_),
    .Y(_03575_));
 AOI21x1_ASAP7_75t_R _09600_ (.A1(_03570_),
    .A2(_03558_),
    .B(_03575_),
    .Y(_03576_));
 NAND2x1_ASAP7_75t_R _09601_ (.A(net3577),
    .B(net3592),
    .Y(_03577_));
 XOR2x2_ASAP7_75t_R _09602_ (.A(_03577_),
    .B(net4078),
    .Y(_03578_));
 NAND2x1_ASAP7_75t_R _09603_ (.A(net3561),
    .B(net3536),
    .Y(_03579_));
 OA21x2_ASAP7_75t_R _09604_ (.A1(net5667),
    .A2(_03578_),
    .B(_03579_),
    .Y(_03580_));
 INVx1_ASAP7_75t_R _09605_ (.A(net3504),
    .Y(_03581_));
 AO21x2_ASAP7_75t_R _09606_ (.A1(net3563),
    .A2(_03560_),
    .B(net5690),
    .Y(_03582_));
 OA31x2_ASAP7_75t_R _09607_ (.A1(net4218),
    .A2(net3632),
    .A3(net3613),
    .B1(net3599),
    .Y(_03583_));
 AOI211x1_ASAP7_75t_R _09608_ (.A1(net3600),
    .A2(net3613),
    .B(net3636),
    .C(net3659),
    .Y(_03584_));
 NOR2x1_ASAP7_75t_R _09609_ (.A(_03583_),
    .B(_03584_),
    .Y(_03585_));
 AO21x1_ASAP7_75t_R _09610_ (.A1(net3550),
    .A2(net3549),
    .B(net3576),
    .Y(_03586_));
 OAI21x1_ASAP7_75t_R _09611_ (.A1(_03582_),
    .A2(net5667),
    .B(_03586_),
    .Y(_03587_));
 XOR2x2_ASAP7_75t_R _09612_ (.A(net3594),
    .B(net3609),
    .Y(_03588_));
 NAND2x1_ASAP7_75t_R _09613_ (.A(_03588_),
    .B(_03585_),
    .Y(_03589_));
 AOI21x1_ASAP7_75t_R _09614_ (.A1(_03560_),
    .A2(net3563),
    .B(_03589_),
    .Y(_03590_));
 XOR2x2_ASAP7_75t_R _09615_ (.A(_03559_),
    .B(_03561_),
    .Y(_03591_));
 NAND2x1_ASAP7_75t_R _09616_ (.A(_03591_),
    .B(net3593),
    .Y(_03592_));
 OAI21x1_ASAP7_75t_R _09617_ (.A1(net3633),
    .A2(net3593),
    .B(_03592_),
    .Y(_03593_));
 XOR2x2_ASAP7_75t_R _09618_ (.A(net3563),
    .B(_03593_),
    .Y(_03594_));
 OAI21x1_ASAP7_75t_R _09619_ (.A1(net3549),
    .A2(_03590_),
    .B(_03594_),
    .Y(_03595_));
 NAND2x1p5_ASAP7_75t_R _09620_ (.A(net3560),
    .B(net5668),
    .Y(_03596_));
 NAND2x2_ASAP7_75t_R _09621_ (.A(_03595_),
    .B(_03596_),
    .Y(_03597_));
 NOR2x2_ASAP7_75t_R _09622_ (.A(_03587_),
    .B(_03597_),
    .Y(_03598_));
 OR3x1_ASAP7_75t_R _09623_ (.A(_03278_),
    .B(net4373),
    .C(net4372),
    .Y(_03599_));
 XNOR2x2_ASAP7_75t_R _09624_ (.A(net4469),
    .B(_03599_),
    .Y(_03600_));
 OAI21x1_ASAP7_75t_R _09625_ (.A1(net3549),
    .A2(_03590_),
    .B(net4078),
    .Y(_03601_));
 NAND2x2_ASAP7_75t_R _09626_ (.A(net4144),
    .B(net5667),
    .Y(_03602_));
 INVx1_ASAP7_75t_R _09627_ (.A(_03577_),
    .Y(_03603_));
 AOI21x1_ASAP7_75t_R _09628_ (.A1(_03602_),
    .A2(_03601_),
    .B(_03603_),
    .Y(_03604_));
 NAND2x2_ASAP7_75t_R _09629_ (.A(net4273),
    .B(_03604_),
    .Y(_03605_));
 NOR2x1_ASAP7_75t_R _09630_ (.A(_03582_),
    .B(net5667),
    .Y(_03606_));
 INVx1_ASAP7_75t_R _09631_ (.A(net3563),
    .Y(_03607_));
 OAI21x1_ASAP7_75t_R _09632_ (.A1(net3633),
    .A2(_03607_),
    .B(net3551),
    .Y(_03608_));
 OA21x2_ASAP7_75t_R _09633_ (.A1(_03606_),
    .A2(net3575),
    .B(_03608_),
    .Y(_03609_));
 AOI21x1_ASAP7_75t_R _09634_ (.A1(_03598_),
    .A2(_03605_),
    .B(_03609_),
    .Y(_03610_));
 NAND2x1_ASAP7_75t_R _09635_ (.A(net5674),
    .B(_03581_),
    .Y(_03611_));
 INVx1_ASAP7_75t_R _09636_ (.A(_03600_),
    .Y(_03612_));
 AOI21x1_ASAP7_75t_R _09637_ (.A1(_03601_),
    .A2(net5984),
    .B(_03612_),
    .Y(_03613_));
 XNOR2x2_ASAP7_75t_R _09638_ (.A(_03613_),
    .B(_03580_),
    .Y(_03614_));
 INVx1_ASAP7_75t_R _09639_ (.A(_03587_),
    .Y(_03615_));
 INVx1_ASAP7_75t_R _09640_ (.A(net5668),
    .Y(_03616_));
 INVx1_ASAP7_75t_R _09641_ (.A(net3560),
    .Y(_03617_));
 AOI211x1_ASAP7_75t_R _09642_ (.A1(net3551),
    .A2(_03607_),
    .B(net3549),
    .C(_03617_),
    .Y(_03618_));
 AOI21x1_ASAP7_75t_R _09643_ (.A1(_03616_),
    .A2(net3548),
    .B(_03618_),
    .Y(_03619_));
 NAND2x1_ASAP7_75t_R _09644_ (.A(_03619_),
    .B(_03615_),
    .Y(_03620_));
 AOI21x1_ASAP7_75t_R _09645_ (.A1(net3562),
    .A2(_03608_),
    .B(net4144),
    .Y(_03621_));
 AOI211x1_ASAP7_75t_R _09646_ (.A1(net3550),
    .A2(net3551),
    .B(net3549),
    .C(net4078),
    .Y(_03622_));
 OAI21x1_ASAP7_75t_R _09647_ (.A1(_03621_),
    .A2(_03622_),
    .B(net3561),
    .Y(_03623_));
 NOR2x1_ASAP7_75t_R _09648_ (.A(_03612_),
    .B(_03623_),
    .Y(_03624_));
 INVx2_ASAP7_75t_R _09649_ (.A(_03609_),
    .Y(_03625_));
 OAI21x1_ASAP7_75t_R _09650_ (.A1(_03624_),
    .A2(_03620_),
    .B(_03625_),
    .Y(_03626_));
 NAND2x1_ASAP7_75t_R _09651_ (.A(_03614_),
    .B(_03626_),
    .Y(_03627_));
 NAND2x1p5_ASAP7_75t_R _09652_ (.A(_03627_),
    .B(_03611_),
    .Y(_03628_));
 AO21x1_ASAP7_75t_R _09653_ (.A1(_03240_),
    .A2(net4468),
    .B(net4276),
    .Y(_03629_));
 XNOR2x2_ASAP7_75t_R _09654_ (.A(net4523),
    .B(_03629_),
    .Y(_03630_));
 INVx1_ASAP7_75t_R _09655_ (.A(_03630_),
    .Y(_03631_));
 AOI211x1_ASAP7_75t_R _09656_ (.A1(net5974),
    .A2(_03623_),
    .B(net3502),
    .C(net4217),
    .Y(_03632_));
 OAI21x1_ASAP7_75t_R _09657_ (.A1(net4217),
    .A2(_03623_),
    .B(net5974),
    .Y(_03633_));
 AOI21x1_ASAP7_75t_R _09658_ (.A1(net3490),
    .A2(_03633_),
    .B(net4273),
    .Y(_03634_));
 NAND2x1_ASAP7_75t_R _09659_ (.A(net3535),
    .B(net3517),
    .Y(_03635_));
 OAI21x1_ASAP7_75t_R _09660_ (.A1(_03632_),
    .A2(_03634_),
    .B(net3499),
    .Y(_03636_));
 NOR2x1_ASAP7_75t_R _09661_ (.A(_03631_),
    .B(_03636_),
    .Y(_03637_));
 NOR2x1_ASAP7_75t_R _09662_ (.A(net3462),
    .B(_03637_),
    .Y(_03638_));
 OAI21x1_ASAP7_75t_R _09663_ (.A1(_03598_),
    .A2(_03609_),
    .B(_03605_),
    .Y(_03639_));
 XOR2x2_ASAP7_75t_R _09664_ (.A(_03639_),
    .B(net3503),
    .Y(_03640_));
 XOR2x2_ASAP7_75t_R _09665_ (.A(_03613_),
    .B(_03580_),
    .Y(_03641_));
 NOR2x1_ASAP7_75t_R _09666_ (.A(_03641_),
    .B(_03610_),
    .Y(_03642_));
 NOR2x1_ASAP7_75t_R _09667_ (.A(_03626_),
    .B(net3504),
    .Y(_03643_));
 NOR2x1_ASAP7_75t_R _09668_ (.A(_03642_),
    .B(_03643_),
    .Y(_03644_));
 NAND2x1_ASAP7_75t_R _09669_ (.A(_03640_),
    .B(_03644_),
    .Y(_03645_));
 NOR2x1_ASAP7_75t_R _09670_ (.A(net3503),
    .B(_03639_),
    .Y(_03646_));
 OA21x2_ASAP7_75t_R _09671_ (.A1(_03646_),
    .A2(net3501),
    .B(net3481),
    .Y(_03647_));
 INVx2_ASAP7_75t_R _09672_ (.A(_03647_),
    .Y(_03648_));
 OAI21x1_ASAP7_75t_R _09673_ (.A1(_03645_),
    .A2(_03637_),
    .B(_03648_),
    .Y(_03649_));
 NAND2x1_ASAP7_75t_R _09674_ (.A(_03638_),
    .B(_03649_),
    .Y(_03650_));
 XOR2x2_ASAP7_75t_R _09675_ (.A(net3473),
    .B(_03650_),
    .Y(_03651_));
 XOR2x2_ASAP7_75t_R _09676_ (.A(_03639_),
    .B(net3500),
    .Y(_03652_));
 NOR2x2_ASAP7_75t_R _09677_ (.A(_03628_),
    .B(_03652_),
    .Y(_03653_));
 NAND2x2_ASAP7_75t_R _09678_ (.A(net4273),
    .B(net5675),
    .Y(_03654_));
 NAND2x1_ASAP7_75t_R _09679_ (.A(net4217),
    .B(_03626_),
    .Y(_03655_));
 INVx1_ASAP7_75t_R _09680_ (.A(net3499),
    .Y(_03656_));
 AOI21x1_ASAP7_75t_R _09681_ (.A1(_03654_),
    .A2(_03655_),
    .B(_03656_),
    .Y(_03657_));
 NAND2x2_ASAP7_75t_R _09682_ (.A(_03657_),
    .B(net4142),
    .Y(_03658_));
 OAI21x1_ASAP7_75t_R _09683_ (.A1(net3458),
    .A2(_03653_),
    .B(_03658_),
    .Y(_03659_));
 XOR2x2_ASAP7_75t_R _09684_ (.A(net3462),
    .B(_03659_),
    .Y(_03660_));
 XOR2x2_ASAP7_75t_R _09685_ (.A(_03635_),
    .B(net4217),
    .Y(_03661_));
 NAND2x2_ASAP7_75t_R _09686_ (.A(_03635_),
    .B(net5675),
    .Y(_03662_));
 OAI21x1_ASAP7_75t_R _09687_ (.A1(_03661_),
    .A2(net3483),
    .B(_03662_),
    .Y(_03663_));
 INVx1_ASAP7_75t_R _09688_ (.A(net3457),
    .Y(_03664_));
 NOR2x2_ASAP7_75t_R _09689_ (.A(_03664_),
    .B(net5701),
    .Y(_03665_));
 OAI21x1_ASAP7_75t_R _09690_ (.A1(net3482),
    .A2(net3474),
    .B(net4142),
    .Y(_03666_));
 XOR2x2_ASAP7_75t_R _09691_ (.A(_03666_),
    .B(_03663_),
    .Y(_03667_));
 AOI21x1_ASAP7_75t_R _09692_ (.A1(_03658_),
    .A2(_03653_),
    .B(_03647_),
    .Y(_03668_));
 NOR2x2_ASAP7_75t_R _09693_ (.A(_03668_),
    .B(_03667_),
    .Y(_03669_));
 NOR2x2_ASAP7_75t_R _09694_ (.A(_03669_),
    .B(_03665_),
    .Y(_03670_));
 NAND2x1p5_ASAP7_75t_R _09695_ (.A(_03660_),
    .B(_03670_),
    .Y(_03671_));
 NAND2x1_ASAP7_75t_R _09696_ (.A(net3472),
    .B(net3471),
    .Y(_03672_));
 INVx1_ASAP7_75t_R _09697_ (.A(_03672_),
    .Y(_03673_));
 AO21x2_ASAP7_75t_R _09698_ (.A1(_03648_),
    .A2(net3443),
    .B(net4142),
    .Y(_03674_));
 INVx2_ASAP7_75t_R _09699_ (.A(_03674_),
    .Y(_03675_));
 AOI211x1_ASAP7_75t_R _09700_ (.A1(net3442),
    .A2(net3461),
    .B(net3459),
    .C(net4077),
    .Y(_03676_));
 NOR2x1_ASAP7_75t_R _09701_ (.A(net4419),
    .B(net4276),
    .Y(_03677_));
 XOR2x2_ASAP7_75t_R _09702_ (.A(_03677_),
    .B(net4465),
    .Y(_03678_));
 OAI21x1_ASAP7_75t_R _09703_ (.A1(_03676_),
    .A2(_03675_),
    .B(_03678_),
    .Y(_03679_));
 NOR2x1p5_ASAP7_75t_R _09704_ (.A(_03673_),
    .B(_03679_),
    .Y(_03680_));
 AOI21x1_ASAP7_75t_R _09705_ (.A1(net3399),
    .A2(net3390),
    .B(net3389),
    .Y(_03681_));
 INVx2_ASAP7_75t_R _09706_ (.A(_03667_),
    .Y(_03682_));
 NAND2x1_ASAP7_75t_R _09707_ (.A(_03682_),
    .B(net3426),
    .Y(_03683_));
 NAND2x1_ASAP7_75t_R _09708_ (.A(net3457),
    .B(_03668_),
    .Y(_03684_));
 NAND2x1_ASAP7_75t_R _09709_ (.A(_03684_),
    .B(_03683_),
    .Y(_03685_));
 XOR2x2_ASAP7_75t_R _09710_ (.A(_03681_),
    .B(net3396),
    .Y(_03686_));
 NOR2x1_ASAP7_75t_R _09711_ (.A(_03673_),
    .B(net3426),
    .Y(_03687_));
 XOR2x2_ASAP7_75t_R _09712_ (.A(_03672_),
    .B(net4077),
    .Y(_03688_));
 NOR2x1_ASAP7_75t_R _09713_ (.A(_03688_),
    .B(net3425),
    .Y(_03689_));
 NOR2x1_ASAP7_75t_R _09714_ (.A(_03687_),
    .B(_03689_),
    .Y(_03690_));
 OAI21x1_ASAP7_75t_R _09715_ (.A1(_03680_),
    .A2(_03671_),
    .B(_03651_),
    .Y(_03691_));
 XOR2x2_ASAP7_75t_R _09716_ (.A(net3397),
    .B(_03690_),
    .Y(_03692_));
 NAND2x1_ASAP7_75t_R _09717_ (.A(_03691_),
    .B(_03692_),
    .Y(_03693_));
 OAI21x1_ASAP7_75t_R _09718_ (.A1(net5676),
    .A2(net3395),
    .B(_03693_),
    .Y(_03694_));
 NAND2x1_ASAP7_75t_R _09719_ (.A(net4143),
    .B(net3424),
    .Y(_03695_));
 NAND2x1_ASAP7_75t_R _09720_ (.A(net3423),
    .B(_03695_),
    .Y(_03696_));
 INVx1_ASAP7_75t_R _09721_ (.A(_03696_),
    .Y(_03697_));
 INVx1_ASAP7_75t_R _09722_ (.A(net4141),
    .Y(_03698_));
 NOR2x2_ASAP7_75t_R _09723_ (.A(net4076),
    .B(_03691_),
    .Y(_03699_));
 XOR2x2_ASAP7_75t_R _09724_ (.A(_03659_),
    .B(net3460),
    .Y(_03700_));
 NOR2x1_ASAP7_75t_R _09725_ (.A(_03685_),
    .B(_03700_),
    .Y(_03701_));
 OAI21x1_ASAP7_75t_R _09726_ (.A1(net3441),
    .A2(net3397),
    .B(_03701_),
    .Y(_03702_));
 AOI21x1_ASAP7_75t_R _09727_ (.A1(net3400),
    .A2(_03702_),
    .B(net4141),
    .Y(_03703_));
 NAND2x1_ASAP7_75t_R _09728_ (.A(net4323),
    .B(net4330),
    .Y(_03704_));
 XOR2x2_ASAP7_75t_R _09729_ (.A(_03704_),
    .B(net4561),
    .Y(_03705_));
 OAI21x1_ASAP7_75t_R _09730_ (.A1(_03703_),
    .A2(_03699_),
    .B(_03705_),
    .Y(_03706_));
 NOR2x1_ASAP7_75t_R _09731_ (.A(net3388),
    .B(net3348),
    .Y(_03707_));
 NOR2x1_ASAP7_75t_R _09732_ (.A(_03694_),
    .B(_03707_),
    .Y(_03708_));
 XOR2x2_ASAP7_75t_R _09733_ (.A(_03681_),
    .B(net3398),
    .Y(_03709_));
 INVx1_ASAP7_75t_R _09734_ (.A(net3395),
    .Y(_03710_));
 NAND3x1_ASAP7_75t_R _09735_ (.A(net3398),
    .B(net3395),
    .C(net3413),
    .Y(_03711_));
 AOI21x1_ASAP7_75t_R _09736_ (.A1(net3399),
    .A2(_03711_),
    .B(net3397),
    .Y(_03712_));
 OR3x1_ASAP7_75t_R _09737_ (.A(net3399),
    .B(net3441),
    .C(net3397),
    .Y(_03713_));
 OAI21x1_ASAP7_75t_R _09738_ (.A1(_03710_),
    .A2(_03712_),
    .B(_03713_),
    .Y(_03714_));
 OAI21x1_ASAP7_75t_R _09739_ (.A1(net3441),
    .A2(net3397),
    .B(net3398),
    .Y(_03715_));
 OAI21x1_ASAP7_75t_R _09740_ (.A1(net5978),
    .A2(_03715_),
    .B(net3411),
    .Y(_03716_));
 NAND2x2_ASAP7_75t_R _09741_ (.A(_03702_),
    .B(_03716_),
    .Y(_03717_));
 INVx2_ASAP7_75t_R _09742_ (.A(_03717_),
    .Y(_03718_));
 AOI21x1_ASAP7_75t_R _09743_ (.A1(_03709_),
    .A2(_03714_),
    .B(_03718_),
    .Y(_03719_));
 NOR2x1_ASAP7_75t_R _09744_ (.A(_03697_),
    .B(_03691_),
    .Y(_03720_));
 XOR2x2_ASAP7_75t_R _09745_ (.A(_03696_),
    .B(_03698_),
    .Y(_03721_));
 AOI21x1_ASAP7_75t_R _09746_ (.A1(net3423),
    .A2(net3412),
    .B(_03698_),
    .Y(_03722_));
 NAND2x1_ASAP7_75t_R _09747_ (.A(net3456),
    .B(_03722_),
    .Y(_03723_));
 INVx1_ASAP7_75t_R _09748_ (.A(net5996),
    .Y(_03724_));
 AOI21x1_ASAP7_75t_R _09749_ (.A1(_03701_),
    .A2(_03723_),
    .B(_03724_),
    .Y(_03725_));
 NOR2x1_ASAP7_75t_R _09750_ (.A(_03721_),
    .B(_03725_),
    .Y(_03726_));
 OAI21x1_ASAP7_75t_R _09751_ (.A1(_03726_),
    .A2(_03720_),
    .B(_03717_),
    .Y(_03727_));
 NOR2x2_ASAP7_75t_R _09752_ (.A(_03706_),
    .B(_03727_),
    .Y(_03728_));
 NOR2x2_ASAP7_75t_R _09753_ (.A(_03719_),
    .B(_03728_),
    .Y(_03729_));
 NAND2x1p5_ASAP7_75t_R _09754_ (.A(_03708_),
    .B(_03729_),
    .Y(_03730_));
 NAND2x1_ASAP7_75t_R _09755_ (.A(net4076),
    .B(_03691_),
    .Y(_03731_));
 NAND2x1_ASAP7_75t_R _09756_ (.A(net4141),
    .B(net3374),
    .Y(_03732_));
 AOI21x1_ASAP7_75t_R _09757_ (.A1(_03731_),
    .A2(_03732_),
    .B(net3388),
    .Y(_03733_));
 AO21x1_ASAP7_75t_R _09758_ (.A1(_03733_),
    .A2(net4216),
    .B(_03694_),
    .Y(_03734_));
 NOR2x1_ASAP7_75t_R _09759_ (.A(net3365),
    .B(_03734_),
    .Y(_03735_));
 AOI21x1_ASAP7_75t_R _09760_ (.A1(net3365),
    .A2(_03730_),
    .B(_03735_),
    .Y(_03736_));
 INVx3_ASAP7_75t_R _09761_ (.A(_03736_),
    .Y(_03737_));
 NAND3x1_ASAP7_75t_R _09762_ (.A(_03733_),
    .B(net4216),
    .C(_03694_),
    .Y(_03738_));
 NAND2x1_ASAP7_75t_R _09763_ (.A(_03738_),
    .B(_03734_),
    .Y(_03739_));
 NOR2x1_ASAP7_75t_R _09764_ (.A(net3347),
    .B(net3364),
    .Y(_03740_));
 AOI21x1_ASAP7_75t_R _09765_ (.A1(_03729_),
    .A2(_03739_),
    .B(_03740_),
    .Y(_03741_));
 NAND2x1_ASAP7_75t_R _09766_ (.A(net3362),
    .B(net3361),
    .Y(_03742_));
 NOR2x1_ASAP7_75t_R _09767_ (.A(_03686_),
    .B(_03694_),
    .Y(_03743_));
 INVx1_ASAP7_75t_R _09768_ (.A(net4216),
    .Y(_03744_));
 OAI21x1_ASAP7_75t_R _09769_ (.A1(_03743_),
    .A2(net3347),
    .B(_03744_),
    .Y(_03745_));
 OAI21x1_ASAP7_75t_R _09770_ (.A1(net5678),
    .A2(net3334),
    .B(net4216),
    .Y(_03746_));
 BUFx3_ASAP7_75t_R place2973 (.A(net5637),
    .Y(net2973));
 NOR2x1_ASAP7_75t_R _09772_ (.A(net4421),
    .B(net4276),
    .Y(_03748_));
 XNOR2x2_ASAP7_75t_R _09773_ (.A(net4562),
    .B(_03748_),
    .Y(_03749_));
 INVx1_ASAP7_75t_R _09774_ (.A(_03749_),
    .Y(_03750_));
 AOI21x1_ASAP7_75t_R _09775_ (.A1(_03745_),
    .A2(_03746_),
    .B(_03750_),
    .Y(_03751_));
 INVx1_ASAP7_75t_R _09776_ (.A(net5671),
    .Y(_03752_));
 OAI21x1_ASAP7_75t_R _09777_ (.A1(net3374),
    .A2(net3387),
    .B(_03752_),
    .Y(_03753_));
 XOR2x2_ASAP7_75t_R _09778_ (.A(_03753_),
    .B(net3348),
    .Y(_03754_));
 OAI21x1_ASAP7_75t_R _09779_ (.A1(net3365),
    .A2(_03694_),
    .B(net3363),
    .Y(_03755_));
 OAI21x1_ASAP7_75t_R _09780_ (.A1(net3349),
    .A2(net3346),
    .B(_03755_),
    .Y(_03756_));
 OAI21x1_ASAP7_75t_R _09781_ (.A1(net3334),
    .A2(net3332),
    .B(net3331),
    .Y(_03757_));
 OAI21x1_ASAP7_75t_R _09782_ (.A1(_03754_),
    .A2(_03756_),
    .B(_03757_),
    .Y(_03758_));
 AOI21x1_ASAP7_75t_R _09783_ (.A1(_03751_),
    .A2(net3345),
    .B(_03758_),
    .Y(_03759_));
 NAND2x1_ASAP7_75t_R _09784_ (.A(_03741_),
    .B(_03759_),
    .Y(_03760_));
 AOI21x1_ASAP7_75t_R _09785_ (.A1(net5686),
    .A2(_03760_),
    .B(net4139),
    .Y(_03761_));
 AOI211x1_ASAP7_75t_R _09786_ (.A1(_03759_),
    .A2(_03741_),
    .B(net3276),
    .C(net4075),
    .Y(_03762_));
 NAND2x1_ASAP7_75t_R _09787_ (.A(net6003),
    .B(net3313),
    .Y(_03763_));
 OAI21x1_ASAP7_75t_R _09788_ (.A1(_03762_),
    .A2(_03761_),
    .B(_03763_),
    .Y(_03764_));
 INVx1_ASAP7_75t_R _09789_ (.A(_03742_),
    .Y(_03765_));
 AOI211x1_ASAP7_75t_R _09790_ (.A1(_03746_),
    .A2(net3314),
    .B(_03765_),
    .C(net4074),
    .Y(_03766_));
 NAND2x1_ASAP7_75t_R _09791_ (.A(net3275),
    .B(_03766_),
    .Y(_03767_));
 INVx1_ASAP7_75t_R _09792_ (.A(net3292),
    .Y(_03768_));
 XOR2x2_ASAP7_75t_R _09793_ (.A(_03742_),
    .B(net4140),
    .Y(_03769_));
 OAI21x1_ASAP7_75t_R _09794_ (.A1(net3335),
    .A2(net3333),
    .B(net3345),
    .Y(_03770_));
 OAI21x1_ASAP7_75t_R _09795_ (.A1(_03769_),
    .A2(net3312),
    .B(_03770_),
    .Y(_03771_));
 NOR2x1_ASAP7_75t_R _09796_ (.A(net3291),
    .B(_03771_),
    .Y(_03772_));
 AOI21x1_ASAP7_75t_R _09797_ (.A1(net3293),
    .A2(_03772_),
    .B(net5672),
    .Y(_03773_));
 OAI21x1_ASAP7_75t_R _09798_ (.A1(net4140),
    .A2(net3335),
    .B(net3330),
    .Y(_03774_));
 OAI21x1_ASAP7_75t_R _09799_ (.A1(net3349),
    .A2(net3312),
    .B(_03774_),
    .Y(_03775_));
 OAI21x1_ASAP7_75t_R _09800_ (.A1(_03768_),
    .A2(_03773_),
    .B(_03775_),
    .Y(_03776_));
 OAI21x1_ASAP7_75t_R _09801_ (.A1(_03737_),
    .A2(_03766_),
    .B(net3291),
    .Y(_03777_));
 OAI21x1_ASAP7_75t_R _09802_ (.A1(_03736_),
    .A2(_03741_),
    .B(_03759_),
    .Y(_03778_));
 NAND2x1p5_ASAP7_75t_R _09803_ (.A(_03777_),
    .B(_03778_),
    .Y(_03779_));
 AOI21x1_ASAP7_75t_R _09804_ (.A1(_03767_),
    .A2(_03776_),
    .B(_03779_),
    .Y(_03780_));
 INVx1_ASAP7_75t_R _09805_ (.A(_03778_),
    .Y(_03781_));
 OA21x2_ASAP7_75t_R _09806_ (.A1(_03781_),
    .A2(net3293),
    .B(net3264),
    .Y(_03782_));
 NAND2x1_ASAP7_75t_R _09807_ (.A(net4425),
    .B(net4330),
    .Y(_03783_));
 XOR2x2_ASAP7_75t_R _09808_ (.A(_03783_),
    .B(net4622),
    .Y(_03784_));
 INVx2_ASAP7_75t_R _09809_ (.A(_03784_),
    .Y(_03785_));
 AOI211x1_ASAP7_75t_R _09810_ (.A1(net5981),
    .A2(_03780_),
    .B(_03782_),
    .C(net4138),
    .Y(_03786_));
 INVx2_ASAP7_75t_R _09811_ (.A(_03782_),
    .Y(_03787_));
 OAI21x1_ASAP7_75t_R _09812_ (.A1(_03785_),
    .A2(net5981),
    .B(_03780_),
    .Y(_03788_));
 AOI21x1_ASAP7_75t_R _09813_ (.A1(_03788_),
    .A2(_03787_),
    .B(net4215),
    .Y(_03789_));
 AOI21x1_ASAP7_75t_R _09814_ (.A1(net3274),
    .A2(net3294),
    .B(net3276),
    .Y(_03790_));
 NAND2x1_ASAP7_75t_R _09815_ (.A(_03790_),
    .B(net4139),
    .Y(_03791_));
 INVx1_ASAP7_75t_R _09816_ (.A(net3291),
    .Y(_03792_));
 NAND2x1_ASAP7_75t_R _09817_ (.A(_03792_),
    .B(_03741_),
    .Y(_03793_));
 OAI21x1_ASAP7_75t_R _09818_ (.A1(_03766_),
    .A2(_03793_),
    .B(net5686),
    .Y(_03794_));
 NAND2x1_ASAP7_75t_R _09819_ (.A(_03794_),
    .B(net4075),
    .Y(_03795_));
 NAND2x1_ASAP7_75t_R _09820_ (.A(net3242),
    .B(net3232),
    .Y(_03796_));
 OAI21x1_ASAP7_75t_R _09821_ (.A1(_03786_),
    .A2(_03789_),
    .B(_03796_),
    .Y(_03797_));
 NOR2x2_ASAP7_75t_R _09822_ (.A(_03186_),
    .B(_03797_),
    .Y(_03798_));
 NAND2x1p5_ASAP7_75t_R _09823_ (.A(_03780_),
    .B(net5981),
    .Y(_03799_));
 AOI21x1_ASAP7_75t_R _09824_ (.A1(_03787_),
    .A2(_03799_),
    .B(net4138),
    .Y(_03800_));
 NOR2x1_ASAP7_75t_R _09825_ (.A(net4075),
    .B(net3262),
    .Y(_03801_));
 XOR2x2_ASAP7_75t_R _09826_ (.A(_03801_),
    .B(net3290),
    .Y(_03802_));
 AOI21x1_ASAP7_75t_R _09827_ (.A1(_03796_),
    .A2(_03800_),
    .B(_03802_),
    .Y(_03803_));
 INVx1_ASAP7_75t_R _09828_ (.A(_03763_),
    .Y(_03804_));
 AOI21x1_ASAP7_75t_R _09829_ (.A1(_03795_),
    .A2(_03791_),
    .B(_03804_),
    .Y(_03805_));
 INVx1_ASAP7_75t_R _09830_ (.A(_03767_),
    .Y(_03806_));
 INVx1_ASAP7_75t_R _09831_ (.A(net3293),
    .Y(_03807_));
 INVx1_ASAP7_75t_R _09832_ (.A(net3349),
    .Y(_03808_));
 AND3x1_ASAP7_75t_R _09833_ (.A(_03808_),
    .B(net3394),
    .C(net3347),
    .Y(_03809_));
 AOI21x1_ASAP7_75t_R _09834_ (.A1(net3329),
    .A2(net3315),
    .B(net3331),
    .Y(_03810_));
 OAI21x1_ASAP7_75t_R _09835_ (.A1(_03809_),
    .A2(_03810_),
    .B(_03775_),
    .Y(_03811_));
 OAI21x1_ASAP7_75t_R _09836_ (.A1(_03807_),
    .A2(_03811_),
    .B(net3265),
    .Y(_03812_));
 AOI21x1_ASAP7_75t_R _09837_ (.A1(net3292),
    .A2(_03812_),
    .B(net3289),
    .Y(_03813_));
 INVx1_ASAP7_75t_R _09838_ (.A(_03779_),
    .Y(_03814_));
 OAI21x1_ASAP7_75t_R _09839_ (.A1(_03806_),
    .A2(_03813_),
    .B(_03814_),
    .Y(_03815_));
 NOR2x1_ASAP7_75t_R _09840_ (.A(_03815_),
    .B(_03805_),
    .Y(_03816_));
 OAI21x1_ASAP7_75t_R _09841_ (.A1(_03816_),
    .A2(_03782_),
    .B(net4215),
    .Y(_03817_));
 NOR2x1p5_ASAP7_75t_R _09842_ (.A(_03817_),
    .B(net3234),
    .Y(_03818_));
 OAI22x1_ASAP7_75t_R _09843_ (.A1(_03785_),
    .A2(net5981),
    .B1(_03780_),
    .B2(_03782_),
    .Y(_03819_));
 NAND2x1_ASAP7_75t_R _09844_ (.A(net3263),
    .B(net3243),
    .Y(_03820_));
 INVx1_ASAP7_75t_R _09845_ (.A(_03820_),
    .Y(_03821_));
 XOR2x2_ASAP7_75t_R _09846_ (.A(_03819_),
    .B(_03821_),
    .Y(_03822_));
 OAI21x1_ASAP7_75t_R _09847_ (.A1(_03803_),
    .A2(_03818_),
    .B(_03822_),
    .Y(_03823_));
 NOR2x1_ASAP7_75t_R _09848_ (.A(net3167),
    .B(net3156),
    .Y(_03824_));
 INVx1_ASAP7_75t_R _09849_ (.A(_03824_),
    .Y(_03825_));
 NOR2x1p5_ASAP7_75t_R _09850_ (.A(_03803_),
    .B(_03818_),
    .Y(_03826_));
 NOR2x1p5_ASAP7_75t_R _09851_ (.A(_03798_),
    .B(_03826_),
    .Y(_03827_));
 NAND2x1_ASAP7_75t_R _09852_ (.A(_03787_),
    .B(_03788_),
    .Y(_03828_));
 NAND2x1_ASAP7_75t_R _09853_ (.A(net4215),
    .B(_03805_),
    .Y(_03829_));
 AND2x2_ASAP7_75t_R _09854_ (.A(_03829_),
    .B(_03820_),
    .Y(_03830_));
 NAND2x1_ASAP7_75t_R _09855_ (.A(_03828_),
    .B(_03830_),
    .Y(_03831_));
 INVx1_ASAP7_75t_R _09856_ (.A(_03788_),
    .Y(_03832_));
 AOI21x1_ASAP7_75t_R _09857_ (.A1(_03831_),
    .A2(net3233),
    .B(_03832_),
    .Y(_03833_));
 AO21x2_ASAP7_75t_R _09858_ (.A1(_03827_),
    .A2(net3166),
    .B(net3189),
    .Y(_03834_));
 NAND2x2_ASAP7_75t_R _09859_ (.A(_03834_),
    .B(_03825_),
    .Y(_03835_));
 INVx1_ASAP7_75t_R _09860_ (.A(_03827_),
    .Y(_03836_));
 NOR2x1_ASAP7_75t_R _09861_ (.A(net5670),
    .B(net3203),
    .Y(_03837_));
 OAI21x1_ASAP7_75t_R _09862_ (.A1(net3217),
    .A2(net3203),
    .B(_03787_),
    .Y(_03838_));
 OAI21x1_ASAP7_75t_R _09863_ (.A1(_03837_),
    .A2(_03838_),
    .B(net4138),
    .Y(_03839_));
 NAND3x1_ASAP7_75t_R _09864_ (.A(net3204),
    .B(net4215),
    .C(net3219),
    .Y(_03840_));
 INVx1_ASAP7_75t_R _09865_ (.A(_03796_),
    .Y(_03841_));
 AOI21x1_ASAP7_75t_R _09866_ (.A1(_03839_),
    .A2(_03840_),
    .B(_03841_),
    .Y(_03842_));
 NAND2x1_ASAP7_75t_R _09867_ (.A(net4278),
    .B(_03842_),
    .Y(_03843_));
 INVx1_ASAP7_75t_R _09868_ (.A(_03802_),
    .Y(_03844_));
 OAI21x1_ASAP7_75t_R _09869_ (.A1(_03841_),
    .A2(_03817_),
    .B(_03844_),
    .Y(_03845_));
 INVx1_ASAP7_75t_R _09870_ (.A(_03818_),
    .Y(_03846_));
 XOR2x2_ASAP7_75t_R _09871_ (.A(net3202),
    .B(net3231),
    .Y(_03847_));
 AOI21x1_ASAP7_75t_R _09872_ (.A1(_03845_),
    .A2(_03846_),
    .B(_03847_),
    .Y(_03848_));
 AOI21x1_ASAP7_75t_R _09873_ (.A1(_03843_),
    .A2(_03848_),
    .B(_03833_),
    .Y(_03849_));
 INVx2_ASAP7_75t_R _09874_ (.A(_03833_),
    .Y(_03850_));
 OAI21x1_ASAP7_75t_R _09875_ (.A1(_03798_),
    .A2(_03850_),
    .B(net3154),
    .Y(_03851_));
 OAI21x1_ASAP7_75t_R _09876_ (.A1(_03849_),
    .A2(_03836_),
    .B(_03851_),
    .Y(_03852_));
 AOI21x1_ASAP7_75t_R _09877_ (.A1(net3126),
    .A2(net3125),
    .B(net3115),
    .Y(_03853_));
 INVx1_ASAP7_75t_R _09878_ (.A(_03853_),
    .Y(_03854_));
 OR3x1_ASAP7_75t_R _09879_ (.A(net4372),
    .B(net4373),
    .C(_03235_),
    .Y(_03855_));
 XOR2x2_ASAP7_75t_R _09880_ (.A(_03855_),
    .B(net4620),
    .Y(_03856_));
 INVx1_ASAP7_75t_R _09881_ (.A(_03856_),
    .Y(_03857_));
 AO21x1_ASAP7_75t_R _09882_ (.A1(net3155),
    .A2(_03850_),
    .B(net4278),
    .Y(_03858_));
 INVx1_ASAP7_75t_R _09883_ (.A(_03858_),
    .Y(_03859_));
 OAI21x1_ASAP7_75t_R _09884_ (.A1(_03823_),
    .A2(_03798_),
    .B(_03850_),
    .Y(_03860_));
 NOR2x1_ASAP7_75t_R _09885_ (.A(net4220),
    .B(_03860_),
    .Y(_03861_));
 NOR2x1_ASAP7_75t_R _09886_ (.A(net3205),
    .B(net3191),
    .Y(_03862_));
 INVx1_ASAP7_75t_R _09887_ (.A(net3180),
    .Y(_03863_));
 OAI21x1_ASAP7_75t_R _09888_ (.A1(_03859_),
    .A2(_03861_),
    .B(_03863_),
    .Y(_03864_));
 NAND2x1p5_ASAP7_75t_R _09889_ (.A(_03860_),
    .B(net3167),
    .Y(_03865_));
 NOR2x1_ASAP7_75t_R _09890_ (.A(net4220),
    .B(_03862_),
    .Y(_03866_));
 INVx1_ASAP7_75t_R _09891_ (.A(_03866_),
    .Y(_03867_));
 XOR2x2_ASAP7_75t_R _09892_ (.A(net3190),
    .B(net3218),
    .Y(_03868_));
 INVx1_ASAP7_75t_R _09893_ (.A(_03868_),
    .Y(_03869_));
 OAI21x1_ASAP7_75t_R _09894_ (.A1(_03867_),
    .A2(_03849_),
    .B(_03869_),
    .Y(_03870_));
 NAND2x1p5_ASAP7_75t_R _09895_ (.A(_03865_),
    .B(_03870_),
    .Y(_03871_));
 OAI21x1_ASAP7_75t_R _09896_ (.A1(_03857_),
    .A2(_03864_),
    .B(_03871_),
    .Y(_03872_));
 AOI21x1_ASAP7_75t_R _09897_ (.A1(net3116),
    .A2(_03854_),
    .B(_03872_),
    .Y(_03873_));
 INVx1_ASAP7_75t_R _09898_ (.A(_03873_),
    .Y(_03874_));
 NAND2x1_ASAP7_75t_R _09899_ (.A(net4278),
    .B(_03849_),
    .Y(_03875_));
 AOI21x1_ASAP7_75t_R _09900_ (.A1(net3141),
    .A2(_03875_),
    .B(net3180),
    .Y(_03876_));
 AOI21x1_ASAP7_75t_R _09901_ (.A1(net3165),
    .A2(net3140),
    .B(net3179),
    .Y(_03877_));
 INVx1_ASAP7_75t_R _09902_ (.A(_03865_),
    .Y(_03878_));
 INVx1_ASAP7_75t_R _09903_ (.A(net3154),
    .Y(_03879_));
 AOI21x1_ASAP7_75t_R _09904_ (.A1(net3166),
    .A2(net3153),
    .B(_03879_),
    .Y(_03880_));
 AOI21x1_ASAP7_75t_R _09905_ (.A1(_03827_),
    .A2(net3140),
    .B(_03880_),
    .Y(_03881_));
 OAI21x1_ASAP7_75t_R _09906_ (.A1(_03877_),
    .A2(_03878_),
    .B(_03881_),
    .Y(_03882_));
 AOI21x1_ASAP7_75t_R _09907_ (.A1(net4272),
    .A2(net3105),
    .B(_03882_),
    .Y(_03883_));
 AO21x2_ASAP7_75t_R _09908_ (.A1(_03874_),
    .A2(net3115),
    .B(_03883_),
    .Y(_03884_));
 OAI21x1_ASAP7_75t_R _09909_ (.A1(_03859_),
    .A2(_03861_),
    .B(_03856_),
    .Y(_03885_));
 NOR2x1_ASAP7_75t_R _09910_ (.A(net3180),
    .B(_03860_),
    .Y(_03886_));
 XOR2x2_ASAP7_75t_R _09911_ (.A(_03862_),
    .B(net4278),
    .Y(_03887_));
 NOR2x1_ASAP7_75t_R _09912_ (.A(_03887_),
    .B(_03849_),
    .Y(_03888_));
 NOR2x1_ASAP7_75t_R _09913_ (.A(_03886_),
    .B(_03888_),
    .Y(_03889_));
 XOR2x2_ASAP7_75t_R _09914_ (.A(_03885_),
    .B(_03889_),
    .Y(_03890_));
 NAND2x1_ASAP7_75t_R _09915_ (.A(net4272),
    .B(_03876_),
    .Y(_03891_));
 AOI21x1_ASAP7_75t_R _09916_ (.A1(_03870_),
    .A2(_03865_),
    .B(_03852_),
    .Y(_03892_));
 INVx3_ASAP7_75t_R _09917_ (.A(_03835_),
    .Y(_03893_));
 AO21x1_ASAP7_75t_R _09918_ (.A1(_03891_),
    .A2(_03892_),
    .B(_03893_),
    .Y(_03894_));
 AOI211x1_ASAP7_75t_R _09919_ (.A1(_03892_),
    .A2(_03885_),
    .B(_03893_),
    .C(_03889_),
    .Y(_03895_));
 AOI21x1_ASAP7_75t_R _09920_ (.A1(_03890_),
    .A2(_03894_),
    .B(_03895_),
    .Y(_03896_));
 OA21x2_ASAP7_75t_R _09921_ (.A1(_03892_),
    .A2(_03893_),
    .B(_03857_),
    .Y(_03897_));
 AOI211x1_ASAP7_75t_R _09922_ (.A1(_03892_),
    .A2(_03864_),
    .B(_03893_),
    .C(_03857_),
    .Y(_03898_));
 NAND2x1_ASAP7_75t_R _09923_ (.A(net3142),
    .B(net3114),
    .Y(_03899_));
 OAI21x1_ASAP7_75t_R _09924_ (.A1(_03897_),
    .A2(_03898_),
    .B(_03899_),
    .Y(_03900_));
 AOI21x1_ASAP7_75t_R _09925_ (.A1(_03893_),
    .A2(_03891_),
    .B(net3106),
    .Y(_03901_));
 NOR2x1_ASAP7_75t_R _09926_ (.A(_03901_),
    .B(_03873_),
    .Y(_03902_));
 NAND3x1_ASAP7_75t_R _09927_ (.A(net3068),
    .B(net5677),
    .C(net3067),
    .Y(_03903_));
 NAND2x1_ASAP7_75t_R _09928_ (.A(net4618),
    .B(net4330),
    .Y(_03904_));
 XOR2x2_ASAP7_75t_R _09929_ (.A(_03904_),
    .B(net4679),
    .Y(_03905_));
 INVx1_ASAP7_75t_R _09930_ (.A(_03905_),
    .Y(_03906_));
 AOI21x1_ASAP7_75t_R _09931_ (.A1(_03884_),
    .A2(_03903_),
    .B(net4137),
    .Y(_03907_));
 AND3x1_ASAP7_75t_R _09932_ (.A(_03882_),
    .B(_03857_),
    .C(net3116),
    .Y(_03908_));
 NAND2x1_ASAP7_75t_R _09933_ (.A(_03864_),
    .B(_03892_),
    .Y(_03909_));
 AOI21x1_ASAP7_75t_R _09934_ (.A1(net3116),
    .A2(_03909_),
    .B(_03857_),
    .Y(_03910_));
 NOR2x1_ASAP7_75t_R _09935_ (.A(_03908_),
    .B(_03910_),
    .Y(_03911_));
 INVx1_ASAP7_75t_R _09936_ (.A(_03911_),
    .Y(_03912_));
 XOR2x2_ASAP7_75t_R _09937_ (.A(net3039),
    .B(net3051),
    .Y(_03913_));
 INVx1_ASAP7_75t_R _09938_ (.A(net3025),
    .Y(_03914_));
 NOR2x2_ASAP7_75t_R _09939_ (.A(_03906_),
    .B(_03900_),
    .Y(_03915_));
 NAND2x2_ASAP7_75t_R _09940_ (.A(_03896_),
    .B(_03902_),
    .Y(_03916_));
 OAI21x1_ASAP7_75t_R _09941_ (.A1(_03916_),
    .A2(_03915_),
    .B(_03884_),
    .Y(_03917_));
 NOR2x2_ASAP7_75t_R _09942_ (.A(net4214),
    .B(_03917_),
    .Y(_03918_));
 OR3x1_ASAP7_75t_R _09943_ (.A(net4372),
    .B(net4373),
    .C(net4676),
    .Y(_03919_));
 XOR2x2_ASAP7_75t_R _09944_ (.A(_03919_),
    .B(net4732),
    .Y(_03920_));
 INVx1_ASAP7_75t_R _09945_ (.A(_03920_),
    .Y(_03921_));
 NOR2x1_ASAP7_75t_R _09946_ (.A(_03921_),
    .B(_03912_),
    .Y(_03922_));
 INVx1_ASAP7_75t_R _09947_ (.A(_03922_),
    .Y(_03923_));
 NOR3x2_ASAP7_75t_R _09948_ (.B(_03907_),
    .C(_03923_),
    .Y(_03924_),
    .A(_03918_));
 INVx3_ASAP7_75t_R _09949_ (.A(_03924_),
    .Y(_03925_));
 AND2x4_ASAP7_75t_R _09950_ (.A(_03917_),
    .B(net3065),
    .Y(_03926_));
 INVx2_ASAP7_75t_R _09951_ (.A(_03926_),
    .Y(_03927_));
 INVx1_ASAP7_75t_R _09952_ (.A(_03884_),
    .Y(_03928_));
 INVx1_ASAP7_75t_R _09953_ (.A(net3067),
    .Y(_03929_));
 OAI21x1_ASAP7_75t_R _09954_ (.A1(net3104),
    .A2(_03883_),
    .B(_03890_),
    .Y(_03930_));
 INVx1_ASAP7_75t_R _09955_ (.A(_03895_),
    .Y(_03931_));
 NAND2x1_ASAP7_75t_R _09956_ (.A(_03930_),
    .B(_03931_),
    .Y(_03932_));
 AOI211x1_ASAP7_75t_R _09957_ (.A1(net3066),
    .A2(net3103),
    .B(_03929_),
    .C(net3063),
    .Y(_03933_));
 OAI21x1_ASAP7_75t_R _09958_ (.A1(_03928_),
    .A2(_03933_),
    .B(net4214),
    .Y(_03934_));
 XOR2x2_ASAP7_75t_R _09959_ (.A(net3079),
    .B(net3103),
    .Y(_03935_));
 INVx1_ASAP7_75t_R _09960_ (.A(_03935_),
    .Y(_03936_));
 OAI21x1_ASAP7_75t_R _09961_ (.A1(net3051),
    .A2(_03934_),
    .B(_03936_),
    .Y(_03937_));
 OA21x2_ASAP7_75t_R _09962_ (.A1(net3064),
    .A2(_03884_),
    .B(_03932_),
    .Y(_03938_));
 INVx1_ASAP7_75t_R _09963_ (.A(_03938_),
    .Y(_03939_));
 NOR2x1_ASAP7_75t_R _09964_ (.A(_03932_),
    .B(net3064),
    .Y(_03940_));
 NAND2x1_ASAP7_75t_R _09965_ (.A(_03940_),
    .B(_03917_),
    .Y(_03941_));
 NAND2x1_ASAP7_75t_R _09966_ (.A(_03939_),
    .B(_03941_),
    .Y(_03942_));
 AOI21x1_ASAP7_75t_R _09967_ (.A1(_03927_),
    .A2(_03937_),
    .B(_03942_),
    .Y(_03943_));
 NOR2x1_ASAP7_75t_R _09968_ (.A(net3065),
    .B(net3050),
    .Y(_03944_));
 AO21x2_ASAP7_75t_R _09969_ (.A1(net3049),
    .A2(_03941_),
    .B(_03944_),
    .Y(_03945_));
 INVx2_ASAP7_75t_R _09970_ (.A(_03945_),
    .Y(_03946_));
 AOI21x1_ASAP7_75t_R _09971_ (.A1(_03925_),
    .A2(_03943_),
    .B(_03946_),
    .Y(_03947_));
 NAND2x1_ASAP7_75t_R _09972_ (.A(_03914_),
    .B(net2995),
    .Y(_03948_));
 NOR2x1_ASAP7_75t_R _09973_ (.A(net4137),
    .B(net3038),
    .Y(_03949_));
 AND2x2_ASAP7_75t_R _09974_ (.A(net3038),
    .B(net4137),
    .Y(_03950_));
 OAI21x1_ASAP7_75t_R _09975_ (.A1(_03949_),
    .A2(_03950_),
    .B(net4271),
    .Y(_03951_));
 XOR2x2_ASAP7_75t_R _09976_ (.A(_03913_),
    .B(_03951_),
    .Y(_03952_));
 AOI21x1_ASAP7_75t_R _09977_ (.A1(net3066),
    .A2(_03907_),
    .B(_03935_),
    .Y(_03953_));
 AOI21x1_ASAP7_75t_R _09978_ (.A1(net3048),
    .A2(_03917_),
    .B(_03938_),
    .Y(_03954_));
 OAI21x1_ASAP7_75t_R _09979_ (.A1(_03926_),
    .A2(_03953_),
    .B(_03954_),
    .Y(_03955_));
 OAI21x1_ASAP7_75t_R _09980_ (.A1(_03924_),
    .A2(_03955_),
    .B(_03945_),
    .Y(_03956_));
 NAND2x1_ASAP7_75t_R _09981_ (.A(_03952_),
    .B(net3002),
    .Y(_03957_));
 AND2x2_ASAP7_75t_R _09982_ (.A(_03948_),
    .B(_03957_),
    .Y(_03958_));
 OAI21x1_ASAP7_75t_R _09983_ (.A1(net3014),
    .A2(net2995),
    .B(net3025),
    .Y(_03959_));
 INVx1_ASAP7_75t_R _09984_ (.A(_03951_),
    .Y(_03960_));
 NAND3x1_ASAP7_75t_R _09985_ (.A(net3001),
    .B(net3066),
    .C(_03960_),
    .Y(_03961_));
 NAND2x1_ASAP7_75t_R _09986_ (.A(_03927_),
    .B(_03937_),
    .Y(_03962_));
 AND2x2_ASAP7_75t_R _09987_ (.A(_03962_),
    .B(_03925_),
    .Y(_03963_));
 AOI21x1_ASAP7_75t_R _09988_ (.A1(net3005),
    .A2(net3003),
    .B(_03962_),
    .Y(_03964_));
 AOI21x1_ASAP7_75t_R _09989_ (.A1(_03963_),
    .A2(_03956_),
    .B(_03964_),
    .Y(_03965_));
 INVx1_ASAP7_75t_R _09990_ (.A(_03965_),
    .Y(_03966_));
 AOI21x1_ASAP7_75t_R _09991_ (.A1(_03959_),
    .A2(_03961_),
    .B(_03966_),
    .Y(_03967_));
 NAND2x1_ASAP7_75t_R _09992_ (.A(net3006),
    .B(net3004),
    .Y(_03968_));
 AO21x1_ASAP7_75t_R _09993_ (.A1(_03963_),
    .A2(net3003),
    .B(net3023),
    .Y(_03969_));
 NAND2x2_ASAP7_75t_R _09994_ (.A(_03968_),
    .B(_03969_),
    .Y(_03970_));
 INVx4_ASAP7_75t_R _09995_ (.A(_03970_),
    .Y(_03971_));
 NAND2x1_ASAP7_75t_R _09996_ (.A(net4730),
    .B(net4330),
    .Y(_03972_));
 XOR2x2_ASAP7_75t_R _09997_ (.A(_03972_),
    .B(net4675),
    .Y(_03973_));
 NAND2x1p5_ASAP7_75t_R _09998_ (.A(net4213),
    .B(_03956_),
    .Y(_03974_));
 NAND2x1p5_ASAP7_75t_R _09999_ (.A(_03947_),
    .B(net4271),
    .Y(_03975_));
 NOR2x1_ASAP7_75t_R _10000_ (.A(net3039),
    .B(net3024),
    .Y(_03976_));
 INVx1_ASAP7_75t_R _10001_ (.A(_03976_),
    .Y(_03977_));
 AOI21x1_ASAP7_75t_R _10002_ (.A1(_03975_),
    .A2(_03974_),
    .B(_03977_),
    .Y(_03978_));
 NAND2x1p5_ASAP7_75t_R _10003_ (.A(_03973_),
    .B(_03978_),
    .Y(_03979_));
 OAI21x1_ASAP7_75t_R _10004_ (.A1(net2949),
    .A2(_03971_),
    .B(net2947),
    .Y(_03980_));
 XNOR2x2_ASAP7_75t_R _10005_ (.A(net2968),
    .B(_03980_),
    .Y(_03981_));
 AO21x1_ASAP7_75t_R _10006_ (.A1(net3002),
    .A2(net4271),
    .B(_03976_),
    .Y(_03982_));
 OA21x2_ASAP7_75t_R _10007_ (.A1(net3014),
    .A2(net2995),
    .B(_03982_),
    .Y(_03983_));
 INVx1_ASAP7_75t_R _10008_ (.A(_03973_),
    .Y(_03984_));
 INVx2_ASAP7_75t_R _10009_ (.A(_03978_),
    .Y(_03985_));
 OAI21x1_ASAP7_75t_R _10010_ (.A1(_03984_),
    .A2(_03985_),
    .B(_03967_),
    .Y(_03986_));
 AO21x1_ASAP7_75t_R _10011_ (.A1(net2979),
    .A2(net2994),
    .B(_03984_),
    .Y(_03987_));
 AOI21x1_ASAP7_75t_R _10012_ (.A1(net2967),
    .A2(_03986_),
    .B(net2965),
    .Y(_03988_));
 OR3x1_ASAP7_75t_R _10013_ (.A(_03985_),
    .B(net4136),
    .C(net2967),
    .Y(_03989_));
 OAI21x1_ASAP7_75t_R _10014_ (.A1(net2978),
    .A2(_03988_),
    .B(_03989_),
    .Y(_03990_));
 NAND2x1_ASAP7_75t_R _10015_ (.A(_03981_),
    .B(_03990_),
    .Y(_03991_));
 INVx1_ASAP7_75t_R _10016_ (.A(_03986_),
    .Y(_03992_));
 AND2x2_ASAP7_75t_R _10017_ (.A(_03979_),
    .B(_03958_),
    .Y(_03993_));
 AOI21x1_ASAP7_75t_R _10018_ (.A1(_03971_),
    .A2(_03993_),
    .B(net2980),
    .Y(_03994_));
 NOR2x1p5_ASAP7_75t_R _10019_ (.A(_03992_),
    .B(_03994_),
    .Y(_03995_));
 INVx2_ASAP7_75t_R _10020_ (.A(_03995_),
    .Y(_03996_));
 OR3x1_ASAP7_75t_R _10021_ (.A(net4372),
    .B(net4373),
    .C(_03232_),
    .Y(_03997_));
 XOR2x2_ASAP7_75t_R _10022_ (.A(_03997_),
    .B(net4754),
    .Y(_03998_));
 INVx1_ASAP7_75t_R _10023_ (.A(_03998_),
    .Y(_03999_));
 AO21x1_ASAP7_75t_R _10024_ (.A1(_03991_),
    .A2(_03996_),
    .B(net4211),
    .Y(_04000_));
 XOR2x2_ASAP7_75t_R _10025_ (.A(_03980_),
    .B(net2968),
    .Y(_04001_));
 AOI21x1_ASAP7_75t_R _10026_ (.A1(_03979_),
    .A2(_03967_),
    .B(_03971_),
    .Y(_04002_));
 XOR2x2_ASAP7_75t_R _10027_ (.A(_03983_),
    .B(_03987_),
    .Y(_04003_));
 NAND2x1_ASAP7_75t_R _10028_ (.A(_04002_),
    .B(_03983_),
    .Y(_04004_));
 OAI21x1_ASAP7_75t_R _10029_ (.A1(net2933),
    .A2(_04003_),
    .B(_04004_),
    .Y(_04005_));
 NOR2x1_ASAP7_75t_R _10030_ (.A(_04001_),
    .B(_04005_),
    .Y(_04006_));
 NAND2x1_ASAP7_75t_R _10031_ (.A(net2994),
    .B(net2979),
    .Y(_04007_));
 NAND3x1_ASAP7_75t_R _10032_ (.A(net2980),
    .B(_03948_),
    .C(_03957_),
    .Y(_04008_));
 NOR2x1_ASAP7_75t_R _10033_ (.A(_03985_),
    .B(_04008_),
    .Y(_04009_));
 OAI21x1_ASAP7_75t_R _10034_ (.A1(net2966),
    .A2(_04008_),
    .B(net2967),
    .Y(_04010_));
 OAI21x1_ASAP7_75t_R _10035_ (.A1(_04009_),
    .A2(_04010_),
    .B(net4136),
    .Y(_04011_));
 NAND2x1_ASAP7_75t_R _10036_ (.A(net4212),
    .B(_04002_),
    .Y(_04012_));
 AOI21x1_ASAP7_75t_R _10037_ (.A1(_04011_),
    .A2(_04012_),
    .B(net4270),
    .Y(_04013_));
 NAND2x1_ASAP7_75t_R _10038_ (.A(net2964),
    .B(_04013_),
    .Y(_04014_));
 AOI21x1_ASAP7_75t_R _10039_ (.A1(_04014_),
    .A2(_04006_),
    .B(net2908),
    .Y(_04015_));
 NAND2x1_ASAP7_75t_R _10040_ (.A(net4211),
    .B(_04015_),
    .Y(_04016_));
 NAND2x1_ASAP7_75t_R _10041_ (.A(net2921),
    .B(net2920),
    .Y(_04017_));
 INVx1_ASAP7_75t_R _10042_ (.A(_04017_),
    .Y(_04018_));
 AOI21x1_ASAP7_75t_R _10043_ (.A1(net2875),
    .A2(_04016_),
    .B(_04018_),
    .Y(_04019_));
 NAND2x1_ASAP7_75t_R _10044_ (.A(net4221),
    .B(_04019_),
    .Y(_04020_));
 INVx1_ASAP7_75t_R _10045_ (.A(_04007_),
    .Y(_04021_));
 AOI211x1_ASAP7_75t_R _10046_ (.A1(net2950),
    .A2(_03985_),
    .B(net2948),
    .C(net4136),
    .Y(_04022_));
 AOI21x1_ASAP7_75t_R _10047_ (.A1(net2967),
    .A2(_03986_),
    .B(net4212),
    .Y(_04023_));
 OAI21x1_ASAP7_75t_R _10048_ (.A1(_04022_),
    .A2(_04023_),
    .B(_03999_),
    .Y(_04024_));
 NOR2x2_ASAP7_75t_R _10049_ (.A(_04021_),
    .B(_04024_),
    .Y(_04025_));
 OAI21x1_ASAP7_75t_R _10050_ (.A1(_04025_),
    .A2(_03991_),
    .B(_03996_),
    .Y(_04026_));
 NAND2x1_ASAP7_75t_R _10051_ (.A(net2884),
    .B(net2874),
    .Y(_04027_));
 XOR2x2_ASAP7_75t_R _10052_ (.A(_04007_),
    .B(net4136),
    .Y(_04028_));
 NAND2x1_ASAP7_75t_R _10053_ (.A(net2964),
    .B(net2934),
    .Y(_04029_));
 OA21x2_ASAP7_75t_R _10054_ (.A1(net2934),
    .A2(_04028_),
    .B(_04029_),
    .Y(_04030_));
 OAI21x1_ASAP7_75t_R _10055_ (.A1(net2904),
    .A2(_04015_),
    .B(net2903),
    .Y(_04031_));
 OAI21x1_ASAP7_75t_R _10056_ (.A1(_03996_),
    .A2(_04025_),
    .B(net2907),
    .Y(_04032_));
 NOR2x1_ASAP7_75t_R _10057_ (.A(_04001_),
    .B(_03995_),
    .Y(_04033_));
 AOI21x1_ASAP7_75t_R _10058_ (.A1(net2964),
    .A2(_04013_),
    .B(_04005_),
    .Y(_04034_));
 OAI21x1_ASAP7_75t_R _10059_ (.A1(net2908),
    .A2(_04033_),
    .B(_04034_),
    .Y(_04035_));
 NAND2x1_ASAP7_75t_R _10060_ (.A(_04032_),
    .B(net2873),
    .Y(_04036_));
 AOI21x1_ASAP7_75t_R _10061_ (.A1(_04027_),
    .A2(_04031_),
    .B(_04036_),
    .Y(_04037_));
 XOR2x2_ASAP7_75t_R _10062_ (.A(net2922),
    .B(_04035_),
    .Y(_04038_));
 AOI21x1_ASAP7_75t_R _10063_ (.A1(_04037_),
    .A2(_04020_),
    .B(net2857),
    .Y(_04039_));
 NOR2x1_ASAP7_75t_R _10064_ (.A(_04020_),
    .B(_04039_),
    .Y(_04040_));
 INVx1_ASAP7_75t_R _10065_ (.A(_03170_),
    .Y(_04041_));
 INVx1_ASAP7_75t_R _10066_ (.A(_04000_),
    .Y(_04042_));
 NOR2x1_ASAP7_75t_R _10067_ (.A(_04026_),
    .B(net4270),
    .Y(_04043_));
 NOR2x2_ASAP7_75t_R _10068_ (.A(_04042_),
    .B(net5687),
    .Y(_04044_));
 NOR2x1_ASAP7_75t_R _10069_ (.A(net4135),
    .B(_04044_),
    .Y(_04045_));
 NOR2x1_ASAP7_75t_R _10070_ (.A(_04015_),
    .B(net2885),
    .Y(_04046_));
 INVx1_ASAP7_75t_R _10071_ (.A(_04030_),
    .Y(_04047_));
 AOI21x1_ASAP7_75t_R _10072_ (.A1(net2906),
    .A2(_04026_),
    .B(_04047_),
    .Y(_04048_));
 INVx1_ASAP7_75t_R _10073_ (.A(_04032_),
    .Y(_04049_));
 OAI21x1_ASAP7_75t_R _10074_ (.A1(net2946),
    .A2(net2904),
    .B(net2909),
    .Y(_04050_));
 AOI21x1_ASAP7_75t_R _10075_ (.A1(net2886),
    .A2(net2922),
    .B(_04050_),
    .Y(_04051_));
 NOR2x1_ASAP7_75t_R _10076_ (.A(_04049_),
    .B(_04051_),
    .Y(_04052_));
 OAI21x1_ASAP7_75t_R _10077_ (.A1(_04048_),
    .A2(_04046_),
    .B(_04052_),
    .Y(_04053_));
 OAI21x1_ASAP7_75t_R _10078_ (.A1(_04042_),
    .A2(_04043_),
    .B(net2905),
    .Y(_04054_));
 NOR2x1_ASAP7_75t_R _10079_ (.A(_04041_),
    .B(_04054_),
    .Y(_04055_));
 INVx2_ASAP7_75t_R _10080_ (.A(_04038_),
    .Y(_04056_));
 OAI21x1_ASAP7_75t_R _10081_ (.A1(_04055_),
    .A2(net2828),
    .B(_04056_),
    .Y(_04057_));
 XOR2x2_ASAP7_75t_R _10082_ (.A(_04017_),
    .B(net4211),
    .Y(_04058_));
 NAND2x1_ASAP7_75t_R _10083_ (.A(_04058_),
    .B(net2874),
    .Y(_04059_));
 OA21x2_ASAP7_75t_R _10084_ (.A1(_04018_),
    .A2(net2874),
    .B(_04059_),
    .Y(_04060_));
 INVx1_ASAP7_75t_R _10085_ (.A(_04060_),
    .Y(_04061_));
 AOI21x1_ASAP7_75t_R _10086_ (.A1(_04045_),
    .A2(_04057_),
    .B(_04061_),
    .Y(_04062_));
 NOR2x1_ASAP7_75t_R _10087_ (.A(net2805),
    .B(net2804),
    .Y(_04063_));
 OR3x1_ASAP7_75t_R _10088_ (.A(net4968),
    .B(net4967),
    .C(net4970),
    .Y(_04064_));
 NAND2x1_ASAP7_75t_R _10089_ (.A(_04064_),
    .B(net4330),
    .Y(_04065_));
 XOR2x2_ASAP7_75t_R _10090_ (.A(_04065_),
    .B(net5175),
    .Y(_04066_));
 AO21x2_ASAP7_75t_R _10091_ (.A1(_04056_),
    .A2(_04053_),
    .B(net4221),
    .Y(_04067_));
 INVx3_ASAP7_75t_R _10092_ (.A(_04067_),
    .Y(_04068_));
 AOI211x1_ASAP7_75t_R _10093_ (.A1(_04037_),
    .A2(net5688),
    .B(net5976),
    .C(net4135),
    .Y(_04069_));
 INVx1_ASAP7_75t_R _10094_ (.A(_04044_),
    .Y(_04070_));
 OAI21x1_ASAP7_75t_R _10095_ (.A1(_04068_),
    .A2(_04069_),
    .B(_04070_),
    .Y(_04071_));
 NOR2x1p5_ASAP7_75t_R _10096_ (.A(_04071_),
    .B(_04066_),
    .Y(_04072_));
 NOR2x1_ASAP7_75t_R _10097_ (.A(_04063_),
    .B(net2780),
    .Y(_04073_));
 NOR2x2_ASAP7_75t_R _10098_ (.A(net2856),
    .B(_04048_),
    .Y(_04074_));
 AOI21x1_ASAP7_75t_R _10099_ (.A1(net4221),
    .A2(net2843),
    .B(_04074_),
    .Y(_04075_));
 INVx1_ASAP7_75t_R _10100_ (.A(_04074_),
    .Y(_04076_));
 AOI21x1_ASAP7_75t_R _10101_ (.A1(net2857),
    .A2(_04020_),
    .B(_04076_),
    .Y(_04077_));
 AOI21x1_ASAP7_75t_R _10102_ (.A1(_04075_),
    .A2(_04057_),
    .B(_04077_),
    .Y(_04078_));
 OAI21x1_ASAP7_75t_R _10103_ (.A1(_04040_),
    .A2(_04062_),
    .B(_04078_),
    .Y(_04079_));
 AND3x1_ASAP7_75t_R _10104_ (.A(net2873),
    .B(net2922),
    .C(_04032_),
    .Y(_04080_));
 OAI21x1_ASAP7_75t_R _10105_ (.A1(_04038_),
    .A2(_04080_),
    .B(_04075_),
    .Y(_04081_));
 AOI21x1_ASAP7_75t_R _10106_ (.A1(net4221),
    .A2(net2843),
    .B(net2828),
    .Y(_04082_));
 AO21x2_ASAP7_75t_R _10107_ (.A1(net2858),
    .A2(_04081_),
    .B(_04082_),
    .Y(_04083_));
 OAI21x1_ASAP7_75t_R _10108_ (.A1(_04079_),
    .A2(_04072_),
    .B(_04083_),
    .Y(_04084_));
 NAND2x1_ASAP7_75t_R _10109_ (.A(_04073_),
    .B(net2763),
    .Y(_04085_));
 XOR2x2_ASAP7_75t_R _10110_ (.A(net2802),
    .B(_04085_),
    .Y(_04086_));
 AOI21x1_ASAP7_75t_R _10111_ (.A1(net2789),
    .A2(net2801),
    .B(net2780),
    .Y(_04087_));
 XOR2x2_ASAP7_75t_R _10112_ (.A(_04087_),
    .B(_04063_),
    .Y(_04088_));
 XOR2x2_ASAP7_75t_R _10113_ (.A(_04044_),
    .B(net4135),
    .Y(_04089_));
 OAI21x1_ASAP7_75t_R _10114_ (.A1(net2857),
    .A2(_04082_),
    .B(_04089_),
    .Y(_04090_));
 OAI21x1_ASAP7_75t_R _10115_ (.A1(net2818),
    .A2(net2842),
    .B(_04090_),
    .Y(_04091_));
 INVx1_ASAP7_75t_R _10116_ (.A(_04066_),
    .Y(_04092_));
 OAI21x1_ASAP7_75t_R _10117_ (.A1(net2803),
    .A2(net2826),
    .B(_04092_),
    .Y(_04093_));
 XOR2x2_ASAP7_75t_R _10118_ (.A(_04091_),
    .B(_04093_),
    .Y(_04094_));
 INVx2_ASAP7_75t_R _10119_ (.A(_04094_),
    .Y(_04095_));
 NAND2x1_ASAP7_75t_R _10120_ (.A(_04084_),
    .B(_04095_),
    .Y(_04096_));
 NAND2x1_ASAP7_75t_R _10121_ (.A(net2827),
    .B(net2817),
    .Y(_04097_));
 INVx1_ASAP7_75t_R _10122_ (.A(net2829),
    .Y(_04098_));
 OAI21x1_ASAP7_75t_R _10123_ (.A1(_04098_),
    .A2(_04039_),
    .B(net2840),
    .Y(_04099_));
 OAI21x1_ASAP7_75t_R _10124_ (.A1(net2841),
    .A2(net2827),
    .B(net2839),
    .Y(_04100_));
 NAND2x1_ASAP7_75t_R _10125_ (.A(_04100_),
    .B(net2815),
    .Y(_04101_));
 AOI21x1_ASAP7_75t_R _10126_ (.A1(_04097_),
    .A2(_04099_),
    .B(_04101_),
    .Y(_04102_));
 INVx1_ASAP7_75t_R _10127_ (.A(net2790),
    .Y(_04103_));
 NAND2x1_ASAP7_75t_R _10128_ (.A(net4134),
    .B(_04103_),
    .Y(_04104_));
 INVx1_ASAP7_75t_R _10129_ (.A(_04083_),
    .Y(_04105_));
 AOI21x1_ASAP7_75t_R _10130_ (.A1(_04102_),
    .A2(_04104_),
    .B(_04105_),
    .Y(_04106_));
 NAND2x1_ASAP7_75t_R _10131_ (.A(net2788),
    .B(_04106_),
    .Y(_04107_));
 NAND2x1_ASAP7_75t_R _10132_ (.A(_04096_),
    .B(_04107_),
    .Y(_04108_));
 NAND2x1_ASAP7_75t_R _10133_ (.A(_04088_),
    .B(_04108_),
    .Y(_04109_));
 NAND2x1_ASAP7_75t_R _10134_ (.A(net4868),
    .B(net4330),
    .Y(_04110_));
 XOR2x2_ASAP7_75t_R _10135_ (.A(_04110_),
    .B(net5176),
    .Y(_04111_));
 INVx1_ASAP7_75t_R _10136_ (.A(_04111_),
    .Y(_04112_));
 AND3x1_ASAP7_75t_R _10137_ (.A(_04112_),
    .B(net5189),
    .C(_00528_),
    .Y(_04113_));
 INVx1_ASAP7_75t_R _10138_ (.A(_04113_),
    .Y(_04114_));
 INVx1_ASAP7_75t_R _10139_ (.A(net2826),
    .Y(_04115_));
 NAND2x1_ASAP7_75t_R _10140_ (.A(net2816),
    .B(_04115_),
    .Y(_04116_));
 INVx1_ASAP7_75t_R _10141_ (.A(_04116_),
    .Y(_04117_));
 NOR2x1_ASAP7_75t_R _10142_ (.A(_04114_),
    .B(_04117_),
    .Y(_04118_));
 INVx1_ASAP7_75t_R _10143_ (.A(_04118_),
    .Y(_04119_));
 XOR2x2_ASAP7_75t_R _10144_ (.A(_04084_),
    .B(net4210),
    .Y(_04120_));
 NOR2x1p5_ASAP7_75t_R _10145_ (.A(_04120_),
    .B(_04119_),
    .Y(_04121_));
 INVx2_ASAP7_75t_R _10146_ (.A(_04121_),
    .Y(_04122_));
 NOR2x1p5_ASAP7_75t_R _10147_ (.A(_04122_),
    .B(_04109_),
    .Y(_04123_));
 AOI21x1_ASAP7_75t_R _10148_ (.A1(_04086_),
    .A2(_04123_),
    .B(net4276),
    .Y(_04124_));
 NAND2x2_ASAP7_75t_R _10149_ (.A(_03165_),
    .B(_04124_),
    .Y(_04125_));
 BUFx3_ASAP7_75t_R place2972 (.A(_02231_),
    .Y(net2972));
 AOI21x1_ASAP7_75t_R _10151_ (.A1(_03164_),
    .A2(net2707),
    .B(net5358),
    .Y(_00744_));
 NAND2x1_ASAP7_75t_R _10152_ (.A(net4975),
    .B(net5030),
    .Y(_04127_));
 AO21x1_ASAP7_75t_R _10153_ (.A1(net2757),
    .A2(_04086_),
    .B(net4276),
    .Y(_04128_));
 XOR2x2_ASAP7_75t_R _10154_ (.A(_04116_),
    .B(net4134),
    .Y(_04129_));
 NAND2x2_ASAP7_75t_R _10155_ (.A(_04129_),
    .B(net2764),
    .Y(_04130_));
 INVx1_ASAP7_75t_R _10156_ (.A(_04130_),
    .Y(_04131_));
 NOR2x1_ASAP7_75t_R _10157_ (.A(net2786),
    .B(net2764),
    .Y(_04132_));
 OAI21x1_ASAP7_75t_R _10158_ (.A1(net4209),
    .A2(net2791),
    .B(net2787),
    .Y(_04133_));
 AOI21x1_ASAP7_75t_R _10159_ (.A1(net2801),
    .A2(_04133_),
    .B(net2779),
    .Y(_04134_));
 INVx1_ASAP7_75t_R _10160_ (.A(net2788),
    .Y(_04135_));
 NOR2x2_ASAP7_75t_R _10161_ (.A(_04135_),
    .B(net2764),
    .Y(_04136_));
 OAI22x1_ASAP7_75t_R _10162_ (.A1(_04131_),
    .A2(_04132_),
    .B1(_04134_),
    .B2(_04136_),
    .Y(_04137_));
 NOR2x1_ASAP7_75t_R _10163_ (.A(_00529_),
    .B(net4208),
    .Y(_04138_));
 INVx1_ASAP7_75t_R _10164_ (.A(_04138_),
    .Y(_04139_));
 NOR2x1p5_ASAP7_75t_R _10165_ (.A(_04139_),
    .B(_04120_),
    .Y(_04140_));
 INVx1_ASAP7_75t_R _10166_ (.A(_04140_),
    .Y(_04141_));
 OAI21x1_ASAP7_75t_R _10167_ (.A1(_04137_),
    .A2(_04141_),
    .B(net4330),
    .Y(_04142_));
 AO21x2_ASAP7_75t_R _10168_ (.A1(_04142_),
    .A2(_04128_),
    .B(net5198),
    .Y(_04143_));
 BUFx3_ASAP7_75t_R place2971 (.A(_02245_),
    .Y(net2971));
 AOI21x1_ASAP7_75t_R _10170_ (.A1(net2723),
    .A2(_04127_),
    .B(net5358),
    .Y(_00745_));
 NAND2x1_ASAP7_75t_R _10171_ (.A(net4976),
    .B(net5030),
    .Y(_04145_));
 AOI21x1_ASAP7_75t_R _10172_ (.A1(net2707),
    .A2(_04145_),
    .B(net5358),
    .Y(_00746_));
 NAND2x1_ASAP7_75t_R _10173_ (.A(net4977),
    .B(net5030),
    .Y(_04146_));
 AOI21x1_ASAP7_75t_R _10174_ (.A1(net2723),
    .A2(_04146_),
    .B(net5358),
    .Y(_00747_));
 NAND2x1_ASAP7_75t_R _10175_ (.A(net4978),
    .B(net5030),
    .Y(_04147_));
 AOI21x1_ASAP7_75t_R _10176_ (.A1(net2707),
    .A2(_04147_),
    .B(net5358),
    .Y(_00748_));
 NAND2x1_ASAP7_75t_R _10177_ (.A(net4979),
    .B(net5030),
    .Y(_04148_));
 AOI21x1_ASAP7_75t_R _10178_ (.A1(net2723),
    .A2(_04148_),
    .B(net5358),
    .Y(_00749_));
 NAND2x1_ASAP7_75t_R _10179_ (.A(net4980),
    .B(net5030),
    .Y(_04149_));
 AOI21x1_ASAP7_75t_R _10180_ (.A1(net2707),
    .A2(_04149_),
    .B(net5358),
    .Y(_00750_));
 NAND2x1_ASAP7_75t_R _10181_ (.A(net4981),
    .B(net5030),
    .Y(_04150_));
 AOI21x1_ASAP7_75t_R _10182_ (.A1(net2723),
    .A2(_04150_),
    .B(net5358),
    .Y(_00751_));
 NAND2x1_ASAP7_75t_R _10183_ (.A(net4982),
    .B(net5031),
    .Y(_04151_));
 AOI21x1_ASAP7_75t_R _10184_ (.A1(net2707),
    .A2(_04151_),
    .B(net5358),
    .Y(_00752_));
 BUFx3_ASAP7_75t_R place2970 (.A(net5421),
    .Y(net2970));
 NAND2x1_ASAP7_75t_R _10186_ (.A(net4983),
    .B(net5031),
    .Y(_04153_));
 BUFx3_ASAP7_75t_R place2969 (.A(_02278_),
    .Y(net2969));
 AOI21x1_ASAP7_75t_R _10188_ (.A1(net2724),
    .A2(_04153_),
    .B(net5358),
    .Y(_00753_));
 OA211x2_ASAP7_75t_R _10189_ (.A1(net5202),
    .A2(net4888),
    .B(net4970),
    .C(net5363),
    .Y(_00754_));
 NAND2x1_ASAP7_75t_R _10190_ (.A(net4984),
    .B(net5030),
    .Y(_04155_));
 AOI21x1_ASAP7_75t_R _10191_ (.A1(net2708),
    .A2(_04155_),
    .B(net5358),
    .Y(_00755_));
 NAND2x1_ASAP7_75t_R _10192_ (.A(net4985),
    .B(net5032),
    .Y(_04156_));
 AOI21x1_ASAP7_75t_R _10193_ (.A1(net2724),
    .A2(_04156_),
    .B(net5358),
    .Y(_00756_));
 NAND2x1_ASAP7_75t_R _10194_ (.A(net4986),
    .B(net5032),
    .Y(_04157_));
 AOI21x1_ASAP7_75t_R _10195_ (.A1(_04157_),
    .A2(net2708),
    .B(net5358),
    .Y(_00757_));
 NAND2x1_ASAP7_75t_R _10196_ (.A(net4987),
    .B(net5032),
    .Y(_04158_));
 AOI21x1_ASAP7_75t_R _10197_ (.A1(net2724),
    .A2(_04158_),
    .B(net5358),
    .Y(_00758_));
 NAND2x1_ASAP7_75t_R _10198_ (.A(net4988),
    .B(net5032),
    .Y(_04159_));
 AOI21x1_ASAP7_75t_R _10199_ (.A1(net2708),
    .A2(_04159_),
    .B(net5358),
    .Y(_00759_));
 NAND2x1_ASAP7_75t_R _10200_ (.A(net4989),
    .B(net5032),
    .Y(_04160_));
 AOI21x1_ASAP7_75t_R _10201_ (.A1(net2724),
    .A2(_04160_),
    .B(net5358),
    .Y(_00760_));
 NAND2x1_ASAP7_75t_R _10202_ (.A(net4990),
    .B(net5032),
    .Y(_04161_));
 AOI21x1_ASAP7_75t_R _10203_ (.A1(_04161_),
    .A2(net2708),
    .B(net5358),
    .Y(_00761_));
 NAND2x1_ASAP7_75t_R _10204_ (.A(net4991),
    .B(net5032),
    .Y(_04162_));
 AOI21x1_ASAP7_75t_R _10205_ (.A1(net2724),
    .A2(_04162_),
    .B(net5358),
    .Y(_00762_));
 NAND2x1_ASAP7_75t_R _10206_ (.A(net4992),
    .B(net5032),
    .Y(_04163_));
 AOI21x1_ASAP7_75t_R _10207_ (.A1(net2708),
    .A2(_04163_),
    .B(net5358),
    .Y(_00763_));
 BUFx3_ASAP7_75t_R place2968 (.A(_03958_),
    .Y(net2968));
 NAND2x1_ASAP7_75t_R _10209_ (.A(net4993),
    .B(net5032),
    .Y(_04165_));
 BUFx3_ASAP7_75t_R place2966 (.A(_03978_),
    .Y(net2966));
 AOI21x1_ASAP7_75t_R _10211_ (.A1(net2724),
    .A2(_04165_),
    .B(net5358),
    .Y(_00764_));
 AO21x1_ASAP7_75t_R _10212_ (.A1(net4330),
    .A2(_00530_),
    .B(net5198),
    .Y(_04167_));
 NAND2x1_ASAP7_75t_R _10213_ (.A(net4968),
    .B(net5029),
    .Y(_04168_));
 AOI211x1_ASAP7_75t_R _10214_ (.A1(_04167_),
    .A2(_04168_),
    .B(net4280),
    .C(net5358),
    .Y(_00765_));
 NAND2x1_ASAP7_75t_R _10215_ (.A(net4994),
    .B(net5032),
    .Y(_04169_));
 AOI21x1_ASAP7_75t_R _10216_ (.A1(net2708),
    .A2(_04169_),
    .B(net5358),
    .Y(_00766_));
 NAND2x1_ASAP7_75t_R _10217_ (.A(net4969),
    .B(net5032),
    .Y(_04170_));
 AOI21x1_ASAP7_75t_R _10218_ (.A1(net2724),
    .A2(_04170_),
    .B(net5358),
    .Y(_00767_));
 INVx2_ASAP7_75t_R _10219_ (.A(net4104),
    .Y(_04171_));
 OR3x1_ASAP7_75t_R _10220_ (.A(_04171_),
    .B(_04112_),
    .C(net4276),
    .Y(_04172_));
 AO21x1_ASAP7_75t_R _10221_ (.A1(net4104),
    .A2(net4330),
    .B(net4208),
    .Y(_04173_));
 AO32x1_ASAP7_75t_R _10222_ (.A1(_04172_),
    .A2(net4888),
    .A3(_04173_),
    .B1(net4967),
    .B2(net5028),
    .Y(_04174_));
 AND2x2_ASAP7_75t_R _10223_ (.A(_04174_),
    .B(net5363),
    .Y(_00768_));
 NAND2x1_ASAP7_75t_R _10224_ (.A(net4966),
    .B(net5029),
    .Y(_04175_));
 AND3x1_ASAP7_75t_R _10225_ (.A(_04120_),
    .B(net4330),
    .C(_04114_),
    .Y(_04176_));
 XOR2x2_ASAP7_75t_R _10226_ (.A(net5725),
    .B(net4134),
    .Y(_04177_));
 OA21x2_ASAP7_75t_R _10227_ (.A1(net4276),
    .A2(_04113_),
    .B(_04177_),
    .Y(_04178_));
 OR3x1_ASAP7_75t_R _10228_ (.A(_04178_),
    .B(net5198),
    .C(_04176_),
    .Y(_04179_));
 AOI21x1_ASAP7_75t_R _10229_ (.A1(_04179_),
    .A2(_04175_),
    .B(net5359),
    .Y(_00769_));
 NAND2x1_ASAP7_75t_R _10230_ (.A(net5709),
    .B(net5029),
    .Y(_04180_));
 NOR2x1_ASAP7_75t_R _10231_ (.A(net2753),
    .B(net2745),
    .Y(_04181_));
 INVx1_ASAP7_75t_R _10232_ (.A(_04181_),
    .Y(_04182_));
 AO21x1_ASAP7_75t_R _10233_ (.A1(_04177_),
    .A2(_04138_),
    .B(net4276),
    .Y(_04183_));
 OAI21x1_ASAP7_75t_R _10234_ (.A1(_04182_),
    .A2(_04183_),
    .B(net4887),
    .Y(_04184_));
 AO21x1_ASAP7_75t_R _10235_ (.A1(_04182_),
    .A2(_04183_),
    .B(_04184_),
    .Y(_04185_));
 AOI21x1_ASAP7_75t_R _10236_ (.A1(_04180_),
    .A2(_04185_),
    .B(net5358),
    .Y(_00770_));
 NAND2x1_ASAP7_75t_R _10237_ (.A(net4964),
    .B(net5029),
    .Y(_04186_));
 AO21x1_ASAP7_75t_R _10238_ (.A1(_04177_),
    .A2(net2778),
    .B(net4276),
    .Y(_04187_));
 OAI21x1_ASAP7_75t_R _10239_ (.A1(net2738),
    .A2(_04187_),
    .B(net4887),
    .Y(_04188_));
 AO21x1_ASAP7_75t_R _10240_ (.A1(net2738),
    .A2(_04187_),
    .B(_04188_),
    .Y(_04189_));
 AOI21x1_ASAP7_75t_R _10241_ (.A1(_04186_),
    .A2(_04189_),
    .B(net5359),
    .Y(_00771_));
 NAND2x1_ASAP7_75t_R _10242_ (.A(net4971),
    .B(net5029),
    .Y(_04190_));
 NAND2x1_ASAP7_75t_R _10243_ (.A(net2757),
    .B(net2732),
    .Y(_04191_));
 XNOR2x2_ASAP7_75t_R _10244_ (.A(net2792),
    .B(net2762),
    .Y(_04192_));
 NAND2x1_ASAP7_75t_R _10245_ (.A(net2800),
    .B(net2755),
    .Y(_04193_));
 AOI22x1_ASAP7_75t_R _10246_ (.A1(net2747),
    .A2(net2756),
    .B1(_04193_),
    .B2(net2754),
    .Y(_04194_));
 AOI21x1_ASAP7_75t_R _10247_ (.A1(net5728),
    .A2(_04194_),
    .B(net4276),
    .Y(_04195_));
 AOI21x1_ASAP7_75t_R _10248_ (.A1(_04195_),
    .A2(net2751),
    .B(net5198),
    .Y(_04196_));
 NAND2x1_ASAP7_75t_R _10249_ (.A(_04196_),
    .B(_04191_),
    .Y(_04197_));
 AOI21x1_ASAP7_75t_R _10250_ (.A1(_04197_),
    .A2(_04190_),
    .B(net5359),
    .Y(_00772_));
 NAND2x1_ASAP7_75t_R _10251_ (.A(net4972),
    .B(net5029),
    .Y(_04198_));
 OAI21x1_ASAP7_75t_R _10252_ (.A1(net4276),
    .A2(_04123_),
    .B(net5719),
    .Y(_04199_));
 INVx1_ASAP7_75t_R _10253_ (.A(_04086_),
    .Y(_04200_));
 NOR2x2_ASAP7_75t_R _10254_ (.A(net2752),
    .B(_04134_),
    .Y(_04201_));
 NOR2x1_ASAP7_75t_R _10255_ (.A(_04192_),
    .B(_04201_),
    .Y(_04202_));
 AOI21x1_ASAP7_75t_R _10256_ (.A1(_04202_),
    .A2(net5983),
    .B(net4276),
    .Y(_04203_));
 AOI21x1_ASAP7_75t_R _10257_ (.A1(_04203_),
    .A2(_04200_),
    .B(net5198),
    .Y(_04204_));
 NAND2x1_ASAP7_75t_R _10258_ (.A(_04199_),
    .B(_04204_),
    .Y(_04205_));
 AOI21x1_ASAP7_75t_R _10259_ (.A1(_04205_),
    .A2(_04198_),
    .B(net5359),
    .Y(_00773_));
 NAND2x1_ASAP7_75t_R _10260_ (.A(net4973),
    .B(net5029),
    .Y(_04206_));
 AOI21x1_ASAP7_75t_R _10261_ (.A1(net2723),
    .A2(_04206_),
    .B(net5358),
    .Y(_00774_));
 AO21x1_ASAP7_75t_R _10262_ (.A1(_01135_),
    .A2(_00334_),
    .B(_01004_),
    .Y(_04207_));
 BUFx3_ASAP7_75t_R place2965 (.A(_03987_),
    .Y(net2965));
 BUFx3_ASAP7_75t_R place2964 (.A(_04007_),
    .Y(net2964));
 NAND2x1_ASAP7_75t_R _10265_ (.A(net5171),
    .B(net5023),
    .Y(_04210_));
 NOR2x1p5_ASAP7_75t_R _10266_ (.A(net4855),
    .B(net5016),
    .Y(_04211_));
 AND2x4_ASAP7_75t_R _10267_ (.A(_04211_),
    .B(net5198),
    .Y(_04212_));
 AOI221x1_ASAP7_75t_R _10268_ (.A1(net5171),
    .A2(net4728),
    .B1(_04210_),
    .B2(net4674),
    .C(_06525_),
    .Y(_00775_));
 INVx6_ASAP7_75t_R _10269_ (.A(_04207_),
    .Y(_04213_));
 AND4x1_ASAP7_75t_R _10270_ (.A(_00993_),
    .B(net5146),
    .C(net5145),
    .D(net4672),
    .Y(_04214_));
 INVx2_ASAP7_75t_R _10271_ (.A(_04214_),
    .Y(_04215_));
 INVx1_ASAP7_75t_R _10272_ (.A(net5170),
    .Y(_04216_));
 AO21x1_ASAP7_75t_R _10273_ (.A1(net5199),
    .A2(net4672),
    .B(net5360),
    .Y(_04217_));
 BUFx3_ASAP7_75t_R place2962 (.A(_05183_),
    .Y(net2962));
 INVx6_ASAP7_75t_R _10275_ (.A(_04217_),
    .Y(_04219_));
 OA21x2_ASAP7_75t_R _10276_ (.A1(_04216_),
    .A2(net4617),
    .B(_04219_),
    .Y(_04220_));
 OA21x2_ASAP7_75t_R _10277_ (.A1(net5170),
    .A2(net4559),
    .B(_04220_),
    .Y(_00776_));
 INVx1_ASAP7_75t_R _10278_ (.A(_00132_),
    .Y(_04221_));
 AND3x1_ASAP7_75t_R _10279_ (.A(_00534_),
    .B(_00535_),
    .C(_00113_),
    .Y(_04222_));
 AND3x4_ASAP7_75t_R _10280_ (.A(_04222_),
    .B(_00109_),
    .C(_00110_),
    .Y(_04223_));
 AND3x1_ASAP7_75t_R _10281_ (.A(_00987_),
    .B(_00105_),
    .C(_00108_),
    .Y(_04224_));
 AND3x4_ASAP7_75t_R _10282_ (.A(_04223_),
    .B(_04213_),
    .C(_04224_),
    .Y(_04225_));
 AND3x1_ASAP7_75t_R _10283_ (.A(net4615),
    .B(net5170),
    .C(net5145),
    .Y(_04226_));
 AOI21x1_ASAP7_75t_R _10284_ (.A1(_04221_),
    .A2(_04226_),
    .B(net4616),
    .Y(_04227_));
 OA21x2_ASAP7_75t_R _10285_ (.A1(_04221_),
    .A2(_04226_),
    .B(_04227_),
    .Y(_00777_));
 INVx1_ASAP7_75t_R _10286_ (.A(net5035),
    .Y(_04228_));
 NOR2x1p5_ASAP7_75t_R _10287_ (.A(_04228_),
    .B(_04215_),
    .Y(_04229_));
 INVx1_ASAP7_75t_R _10288_ (.A(_04229_),
    .Y(_04230_));
 INVx1_ASAP7_75t_R _10289_ (.A(net5169),
    .Y(_04231_));
 OA21x2_ASAP7_75t_R _10290_ (.A1(_04231_),
    .A2(_04229_),
    .B(_04219_),
    .Y(_04232_));
 OA21x2_ASAP7_75t_R _10291_ (.A1(net5169),
    .A2(_04230_),
    .B(_04232_),
    .Y(_00778_));
 AND3x1_ASAP7_75t_R _10292_ (.A(_00985_),
    .B(_00131_),
    .C(_00337_),
    .Y(_04233_));
 INVx1_ASAP7_75t_R _10293_ (.A(_04233_),
    .Y(_04234_));
 INVx4_ASAP7_75t_R _10294_ (.A(_04225_),
    .Y(_04235_));
 NOR2x1p5_ASAP7_75t_R _10295_ (.A(net4726),
    .B(net4557),
    .Y(_04236_));
 INVx2_ASAP7_75t_R _10296_ (.A(_04236_),
    .Y(_04237_));
 INVx1_ASAP7_75t_R _10297_ (.A(net5168),
    .Y(_04238_));
 OA21x2_ASAP7_75t_R _10298_ (.A1(net4883),
    .A2(_04236_),
    .B(_04219_),
    .Y(_04239_));
 OA21x2_ASAP7_75t_R _10299_ (.A1(net5168),
    .A2(_04237_),
    .B(_04239_),
    .Y(_00779_));
 OR5x1_ASAP7_75t_R _10300_ (.A(net5167),
    .B(net4559),
    .C(_04238_),
    .D(_04231_),
    .E(_04228_),
    .Y(_04240_));
 BUFx3_ASAP7_75t_R place2961 (.A(_05206_),
    .Y(net2961));
 AND3x1_ASAP7_75t_R _10302_ (.A(net5035),
    .B(net5168),
    .C(net5169),
    .Y(_04242_));
 INVx1_ASAP7_75t_R _10303_ (.A(net5167),
    .Y(_04243_));
 AO21x1_ASAP7_75t_R _10304_ (.A1(net4617),
    .A2(_04242_),
    .B(_04243_),
    .Y(_04244_));
 AND3x1_ASAP7_75t_R _10305_ (.A(_04240_),
    .B(_04219_),
    .C(_04244_),
    .Y(_00780_));
 INVx1_ASAP7_75t_R _10306_ (.A(_00128_),
    .Y(_04245_));
 AND3x1_ASAP7_75t_R _10307_ (.A(_04236_),
    .B(net5167),
    .C(net5168),
    .Y(_04246_));
 OAI21x1_ASAP7_75t_R _10308_ (.A1(_04246_),
    .A2(_04245_),
    .B(_04219_),
    .Y(_04247_));
 AOI21x1_ASAP7_75t_R _10309_ (.A1(_04245_),
    .A2(net4464),
    .B(_04247_),
    .Y(_00781_));
 AND3x1_ASAP7_75t_R _10310_ (.A(net4748),
    .B(net4672),
    .C(net4697),
    .Y(_04248_));
 INVx1_ASAP7_75t_R _10311_ (.A(_04248_),
    .Y(_04249_));
 AOI21x1_ASAP7_75t_R _10312_ (.A1(net5166),
    .A2(_04249_),
    .B(net4616),
    .Y(_04250_));
 OA21x2_ASAP7_75t_R _10313_ (.A1(net5166),
    .A2(net4556),
    .B(_04250_),
    .Y(_00782_));
 AND3x1_ASAP7_75t_R _10314_ (.A(_00983_),
    .B(_00127_),
    .C(_00130_),
    .Y(_04251_));
 INVx1_ASAP7_75t_R _10315_ (.A(_04251_),
    .Y(_04252_));
 OR3x1_ASAP7_75t_R _10316_ (.A(_04237_),
    .B(_00126_),
    .C(net4725),
    .Y(_04253_));
 OAI21x1_ASAP7_75t_R _10317_ (.A1(net4725),
    .A2(_04237_),
    .B(_00126_),
    .Y(_04254_));
 AND3x1_ASAP7_75t_R _10318_ (.A(_04254_),
    .B(_04219_),
    .C(_04253_),
    .Y(_00783_));
 AND3x1_ASAP7_75t_R _10319_ (.A(_04229_),
    .B(_00976_),
    .C(net4858),
    .Y(_04255_));
 INVx1_ASAP7_75t_R _10320_ (.A(_04255_),
    .Y(_04256_));
 OAI21x1_ASAP7_75t_R _10321_ (.A1(net5165),
    .A2(_04256_),
    .B(_04219_),
    .Y(_04257_));
 AOI21x1_ASAP7_75t_R _10322_ (.A1(net5165),
    .A2(_04256_),
    .B(_04257_),
    .Y(_00784_));
 AND2x2_ASAP7_75t_R _10323_ (.A(_00125_),
    .B(_00126_),
    .Y(_04258_));
 INVx1_ASAP7_75t_R _10324_ (.A(_04258_),
    .Y(_04259_));
 OR4x1_ASAP7_75t_R _10325_ (.A(_04235_),
    .B(_04234_),
    .C(_04252_),
    .D(_04259_),
    .Y(_04260_));
 INVx1_ASAP7_75t_R _10326_ (.A(net5164),
    .Y(_04261_));
 AND2x2_ASAP7_75t_R _10327_ (.A(_04260_),
    .B(_04261_),
    .Y(_04262_));
 NOR2x1_ASAP7_75t_R _10328_ (.A(_04261_),
    .B(_04260_),
    .Y(_04263_));
 OA21x2_ASAP7_75t_R _10329_ (.A1(_04262_),
    .A2(_04263_),
    .B(net4558),
    .Y(_00785_));
 NAND2x1_ASAP7_75t_R _10330_ (.A(_00537_),
    .B(net5023),
    .Y(_04264_));
 AOI221x1_ASAP7_75t_R _10331_ (.A1(net5163),
    .A2(net4728),
    .B1(_04264_),
    .B2(net4674),
    .C(_06525_),
    .Y(_00786_));
 AND3x1_ASAP7_75t_R _10332_ (.A(_04229_),
    .B(_00977_),
    .C(net4858),
    .Y(_04265_));
 INVx2_ASAP7_75t_R _10333_ (.A(net4463),
    .Y(_04266_));
 AOI21x1_ASAP7_75t_R _10334_ (.A1(net5162),
    .A2(_04266_),
    .B(net4616),
    .Y(_04267_));
 OA21x2_ASAP7_75t_R _10335_ (.A1(net5162),
    .A2(_04266_),
    .B(_04267_),
    .Y(_00787_));
 AND4x1_ASAP7_75t_R _10336_ (.A(net4839),
    .B(net5162),
    .C(net5164),
    .D(_04258_),
    .Y(_04268_));
 AND3x1_ASAP7_75t_R _10337_ (.A(_04268_),
    .B(_04233_),
    .C(net4615),
    .Y(_04269_));
 INVx1_ASAP7_75t_R _10338_ (.A(_04269_),
    .Y(_04270_));
 INVx1_ASAP7_75t_R _10339_ (.A(net5161),
    .Y(_04271_));
 OA21x2_ASAP7_75t_R _10340_ (.A1(_04271_),
    .A2(_04269_),
    .B(_04219_),
    .Y(_04272_));
 OA21x2_ASAP7_75t_R _10341_ (.A1(net5161),
    .A2(_04270_),
    .B(_04272_),
    .Y(_00788_));
 AND3x1_ASAP7_75t_R _10342_ (.A(_04265_),
    .B(net5161),
    .C(net5162),
    .Y(_04273_));
 INVx1_ASAP7_75t_R _10343_ (.A(_04273_),
    .Y(_04274_));
 INVx1_ASAP7_75t_R _10344_ (.A(net5160),
    .Y(_04275_));
 OA21x2_ASAP7_75t_R _10345_ (.A1(_04275_),
    .A2(_04273_),
    .B(_04219_),
    .Y(_04276_));
 OA21x2_ASAP7_75t_R _10346_ (.A1(_04274_),
    .A2(net5160),
    .B(_04276_),
    .Y(_00789_));
 AND3x1_ASAP7_75t_R _10347_ (.A(_04263_),
    .B(net5160),
    .C(_00974_),
    .Y(_04277_));
 XOR2x2_ASAP7_75t_R _10348_ (.A(net4417),
    .B(net5159),
    .Y(_04278_));
 NOR2x1_ASAP7_75t_R _10349_ (.A(net4616),
    .B(_04278_),
    .Y(_00790_));
 INVx1_ASAP7_75t_R _10350_ (.A(net4749),
    .Y(_04279_));
 OR3x1_ASAP7_75t_R _10351_ (.A(_04249_),
    .B(_00119_),
    .C(_04279_),
    .Y(_04280_));
 INVx1_ASAP7_75t_R _10352_ (.A(_00119_),
    .Y(_04281_));
 AO21x1_ASAP7_75t_R _10353_ (.A1(_04248_),
    .A2(net4749),
    .B(_04281_),
    .Y(_04282_));
 AND3x1_ASAP7_75t_R _10354_ (.A(_04280_),
    .B(_04219_),
    .C(_04282_),
    .Y(_00791_));
 AND3x1_ASAP7_75t_R _10355_ (.A(_04277_),
    .B(_00119_),
    .C(net5159),
    .Y(_04283_));
 XOR2x2_ASAP7_75t_R _10356_ (.A(net4364),
    .B(net5158),
    .Y(_04284_));
 NOR2x1_ASAP7_75t_R _10357_ (.A(net4616),
    .B(_04284_),
    .Y(_00792_));
 AND3x1_ASAP7_75t_R _10358_ (.A(_00979_),
    .B(net5159),
    .C(net5160),
    .Y(_04285_));
 INVx1_ASAP7_75t_R _10359_ (.A(_04285_),
    .Y(_04286_));
 NOR2x1_ASAP7_75t_R _10360_ (.A(_04286_),
    .B(_04274_),
    .Y(_04287_));
 INVx2_ASAP7_75t_R _10361_ (.A(_04287_),
    .Y(_04288_));
 OAI21x1_ASAP7_75t_R _10362_ (.A1(net5157),
    .A2(net4269),
    .B(_04219_),
    .Y(_04289_));
 AOI21x1_ASAP7_75t_R _10363_ (.A1(net5157),
    .A2(net4269),
    .B(_04289_),
    .Y(_00793_));
 AND3x1_ASAP7_75t_R _10364_ (.A(_04283_),
    .B(net5157),
    .C(net5158),
    .Y(_04290_));
 XOR2x2_ASAP7_75t_R _10365_ (.A(net4322),
    .B(net5156),
    .Y(_04291_));
 NOR2x1_ASAP7_75t_R _10366_ (.A(net4616),
    .B(_04291_),
    .Y(_00794_));
 AND2x2_ASAP7_75t_R _10367_ (.A(net4859),
    .B(_00980_),
    .Y(_04292_));
 INVx1_ASAP7_75t_R _10368_ (.A(_04292_),
    .Y(_04293_));
 OR3x1_ASAP7_75t_R _10369_ (.A(_04266_),
    .B(net5155),
    .C(_04293_),
    .Y(_04294_));
 OAI21x1_ASAP7_75t_R _10370_ (.A1(_04293_),
    .A2(_04266_),
    .B(net5155),
    .Y(_04295_));
 AND3x1_ASAP7_75t_R _10371_ (.A(_04295_),
    .B(_04219_),
    .C(_04294_),
    .Y(_00795_));
 INVx1_ASAP7_75t_R _10372_ (.A(net5154),
    .Y(_04296_));
 AND3x1_ASAP7_75t_R _10373_ (.A(_04290_),
    .B(net5155),
    .C(net5156),
    .Y(_04297_));
 INVx1_ASAP7_75t_R _10374_ (.A(_04297_),
    .Y(_04298_));
 OA21x2_ASAP7_75t_R _10375_ (.A1(_04298_),
    .A2(net5154),
    .B(_04219_),
    .Y(_04299_));
 OA21x2_ASAP7_75t_R _10376_ (.A1(_04296_),
    .A2(_04297_),
    .B(_04299_),
    .Y(_00796_));
 OAI21x1_ASAP7_75t_R _10377_ (.A1(net4867),
    .A2(net5153),
    .B(net5023),
    .Y(_04300_));
 AO21x1_ASAP7_75t_R _10378_ (.A1(_04212_),
    .A2(net4867),
    .B(net4728),
    .Y(_04301_));
 AOI221x1_ASAP7_75t_R _10379_ (.A1(net4673),
    .A2(_04300_),
    .B1(net5153),
    .B2(_04301_),
    .C(_06525_),
    .Y(_00797_));
 AND4x1_ASAP7_75t_R _10380_ (.A(net5154),
    .B(net5155),
    .C(net5156),
    .D(net5157),
    .Y(_04302_));
 INVx1_ASAP7_75t_R _10381_ (.A(_04302_),
    .Y(_04303_));
 OR3x1_ASAP7_75t_R _10382_ (.A(_04288_),
    .B(net5152),
    .C(_04303_),
    .Y(_04304_));
 OAI21x1_ASAP7_75t_R _10383_ (.A1(_04303_),
    .A2(_04288_),
    .B(net5152),
    .Y(_04305_));
 AND3x1_ASAP7_75t_R _10384_ (.A(_04304_),
    .B(_04219_),
    .C(_04305_),
    .Y(_00798_));
 INVx1_ASAP7_75t_R _10385_ (.A(_00981_),
    .Y(_04306_));
 OR3x1_ASAP7_75t_R _10386_ (.A(_04298_),
    .B(_00111_),
    .C(_04306_),
    .Y(_04307_));
 OAI21x1_ASAP7_75t_R _10387_ (.A1(_04306_),
    .A2(_04298_),
    .B(_00111_),
    .Y(_04308_));
 AND3x1_ASAP7_75t_R _10388_ (.A(_04307_),
    .B(_04219_),
    .C(_04308_),
    .Y(_00799_));
 XOR2x2_ASAP7_75t_R _10389_ (.A(net4884),
    .B(net5151),
    .Y(_04309_));
 OAI21x1_ASAP7_75t_R _10390_ (.A1(net5199),
    .A2(_04309_),
    .B(_04212_),
    .Y(_04310_));
 OA211x2_ASAP7_75t_R _10391_ (.A1(_00989_),
    .A2(net4672),
    .B(_04310_),
    .C(net5363),
    .Y(_00800_));
 XNOR2x2_ASAP7_75t_R _10392_ (.A(net5150),
    .B(net4856),
    .Y(_04311_));
 OA21x2_ASAP7_75t_R _10393_ (.A1(_04311_),
    .A2(net5199),
    .B(net5198),
    .Y(_04312_));
 NOR2x1_ASAP7_75t_R _10394_ (.A(net4728),
    .B(_04312_),
    .Y(_04313_));
 NOR2x1_ASAP7_75t_R _10395_ (.A(net5150),
    .B(net4672),
    .Y(_04314_));
 OA21x2_ASAP7_75t_R _10396_ (.A1(_04313_),
    .A2(_04314_),
    .B(net5363),
    .Y(_00801_));
 AND3x1_ASAP7_75t_R _10397_ (.A(net4840),
    .B(net4672),
    .C(net5149),
    .Y(_04315_));
 AOI21x1_ASAP7_75t_R _10398_ (.A1(net4672),
    .A2(net4840),
    .B(net5149),
    .Y(_04316_));
 OA21x2_ASAP7_75t_R _10399_ (.A1(_04315_),
    .A2(_04316_),
    .B(_04219_),
    .Y(_00802_));
 AND3x1_ASAP7_75t_R _10400_ (.A(_00992_),
    .B(net5149),
    .C(net5150),
    .Y(_04317_));
 INVx1_ASAP7_75t_R _10401_ (.A(_04317_),
    .Y(_04318_));
 OR3x1_ASAP7_75t_R _10402_ (.A(_04318_),
    .B(net5148),
    .C(net4728),
    .Y(_04319_));
 OAI21x1_ASAP7_75t_R _10403_ (.A1(net4728),
    .A2(_04318_),
    .B(net5148),
    .Y(_04320_));
 AND3x1_ASAP7_75t_R _10404_ (.A(_04219_),
    .B(_04319_),
    .C(_04320_),
    .Y(_00803_));
 AND3x1_ASAP7_75t_R _10405_ (.A(net4840),
    .B(net5148),
    .C(net5149),
    .Y(_04321_));
 INVx1_ASAP7_75t_R _10406_ (.A(net5147),
    .Y(_04322_));
 AND2x2_ASAP7_75t_R _10407_ (.A(_04321_),
    .B(_04322_),
    .Y(_04323_));
 NOR2x1_ASAP7_75t_R _10408_ (.A(_04322_),
    .B(_04321_),
    .Y(_04324_));
 OR3x1_ASAP7_75t_R _10409_ (.A(_04324_),
    .B(net5200),
    .C(_04323_),
    .Y(_04325_));
 AOI221x1_ASAP7_75t_R _10410_ (.A1(net5147),
    .A2(net4728),
    .B1(net4673),
    .B2(_04325_),
    .C(_06525_),
    .Y(_00804_));
 XOR2x2_ASAP7_75t_R _10411_ (.A(net5146),
    .B(net4697),
    .Y(_04326_));
 OA21x2_ASAP7_75t_R _10412_ (.A1(_04326_),
    .A2(net5200),
    .B(net4727),
    .Y(_04327_));
 AOI211x1_ASAP7_75t_R _10413_ (.A1(net5146),
    .A2(net4728),
    .B(_04327_),
    .C(net5360),
    .Y(_00805_));
 AOI21x1_ASAP7_75t_R _10414_ (.A1(net5145),
    .A2(net4557),
    .B(net4616),
    .Y(_04328_));
 OA21x2_ASAP7_75t_R _10415_ (.A1(net5145),
    .A2(net4557),
    .B(_04328_),
    .Y(_00806_));
 NOR2x2_ASAP7_75t_R _10416_ (.A(_02522_),
    .B(_00175_),
    .Y(_04329_));
 INVx8_ASAP7_75t_R _10417_ (.A(net5504),
    .Y(_04330_));
 BUFx3_ASAP7_75t_R place2960 (.A(_05207_),
    .Y(net2960));
 BUFx3_ASAP7_75t_R place2959 (.A(_06273_),
    .Y(net2959));
 AO21x1_ASAP7_75t_R _10420_ (.A1(net5019),
    .A2(net2710),
    .B(net5359),
    .Y(_04333_));
 AOI21x1_ASAP7_75t_R _10421_ (.A1(net5923),
    .A2(net5143),
    .B(_04333_),
    .Y(_00807_));
 BUFx3_ASAP7_75t_R place2956 (.A(_06346_),
    .Y(net2956));
 NAND2x1_ASAP7_75t_R _10423_ (.A(net4944),
    .B(net2700),
    .Y(_04335_));
 AND3x1_ASAP7_75t_R _10424_ (.A(net5019),
    .B(net4936),
    .C(net4935),
    .Y(_04336_));
 XOR2x2_ASAP7_75t_R _10425_ (.A(net4838),
    .B(net4937),
    .Y(_04337_));
 INVx1_ASAP7_75t_R _10426_ (.A(_04337_),
    .Y(_04338_));
 OR3x1_ASAP7_75t_R _10427_ (.A(_00539_),
    .B(_00079_),
    .C(net5124),
    .Y(_04339_));
 XOR2x2_ASAP7_75t_R _10428_ (.A(net4724),
    .B(net5122),
    .Y(_04340_));
 INVx1_ASAP7_75t_R _10429_ (.A(_04340_),
    .Y(_04341_));
 XOR2x2_ASAP7_75t_R _10430_ (.A(net4816),
    .B(net5124),
    .Y(_04342_));
 INVx1_ASAP7_75t_R _10431_ (.A(_04342_),
    .Y(_04343_));
 AND3x1_ASAP7_75t_R _10432_ (.A(_04343_),
    .B(net5019),
    .C(_00540_),
    .Y(_04344_));
 AND3x1_ASAP7_75t_R _10433_ (.A(net4671),
    .B(net4614),
    .C(_04344_),
    .Y(_04345_));
 INVx1_ASAP7_75t_R _10434_ (.A(net4555),
    .Y(_04346_));
 INVx1_ASAP7_75t_R _10435_ (.A(net5123),
    .Y(_04347_));
 AND4x1_ASAP7_75t_R _10436_ (.A(net4942),
    .B(net4941),
    .C(net4940),
    .D(net4939),
    .Y(_04348_));
 AND3x2_ASAP7_75t_R _10437_ (.A(_04336_),
    .B(net4938),
    .C(net4937),
    .Y(_04349_));
 NAND2x2_ASAP7_75t_R _10438_ (.A(_04348_),
    .B(_04349_),
    .Y(_04350_));
 OR4x1_ASAP7_75t_R _10439_ (.A(net5139),
    .B(net5140),
    .C(net5141),
    .D(net5142),
    .Y(_04351_));
 OR4x1_ASAP7_75t_R _10440_ (.A(_04350_),
    .B(net5117),
    .C(net5138),
    .D(_04351_),
    .Y(_04352_));
 OR3x1_ASAP7_75t_R _10441_ (.A(net5134),
    .B(net5135),
    .C(net5136),
    .Y(_04353_));
 OR4x1_ASAP7_75t_R _10442_ (.A(net5129),
    .B(net5130),
    .C(net5131),
    .D(net5133),
    .Y(_04354_));
 OR4x1_ASAP7_75t_R _10443_ (.A(_04352_),
    .B(net5137),
    .C(_04353_),
    .D(_04354_),
    .Y(_04355_));
 INVx1_ASAP7_75t_R _10444_ (.A(_04355_),
    .Y(_04356_));
 AND3x1_ASAP7_75t_R _10445_ (.A(net4961),
    .B(net4960),
    .C(net4959),
    .Y(_04357_));
 AND3x1_ASAP7_75t_R _10446_ (.A(_04357_),
    .B(net4962),
    .C(net4958),
    .Y(_04358_));
 NOR2x1_ASAP7_75t_R _10447_ (.A(net5127),
    .B(net5128),
    .Y(_04359_));
 AND4x1_ASAP7_75t_R _10448_ (.A(net4518),
    .B(net4963),
    .C(_04358_),
    .D(net4880),
    .Y(_04360_));
 NOR2x1_ASAP7_75t_R _10449_ (.A(_04347_),
    .B(_04360_),
    .Y(_04361_));
 AND2x2_ASAP7_75t_R _10450_ (.A(_04360_),
    .B(_04347_),
    .Y(_04362_));
 NOR2x1_ASAP7_75t_R _10451_ (.A(_04361_),
    .B(_04362_),
    .Y(_04363_));
 BUFx3_ASAP7_75t_R place2955 (.A(_02232_),
    .Y(net2955));
 NAND2x1_ASAP7_75t_R _10453_ (.A(_04346_),
    .B(net4362),
    .Y(_04365_));
 XOR2x2_ASAP7_75t_R _10454_ (.A(net4723),
    .B(net4939),
    .Y(_04366_));
 XOR2x2_ASAP7_75t_R _10455_ (.A(_04365_),
    .B(net4668),
    .Y(_04367_));
 INVx1_ASAP7_75t_R _10456_ (.A(_04367_),
    .Y(_04368_));
 OR3x1_ASAP7_75t_R _10457_ (.A(_04339_),
    .B(net5121),
    .C(net5122),
    .Y(_04369_));
 OR5x1_ASAP7_75t_R _10458_ (.A(net5117),
    .B(net4667),
    .C(net5118),
    .D(net5119),
    .E(net5120),
    .Y(_04370_));
 XOR2x2_ASAP7_75t_R _10459_ (.A(_04370_),
    .B(net5142),
    .Y(_04371_));
 INVx1_ASAP7_75t_R _10460_ (.A(_04371_),
    .Y(_04372_));
 INVx1_ASAP7_75t_R _10461_ (.A(_04369_),
    .Y(_04373_));
 AND3x1_ASAP7_75t_R _10462_ (.A(_04373_),
    .B(net4941),
    .C(net4940),
    .Y(_04374_));
 XOR2x2_ASAP7_75t_R _10463_ (.A(_04374_),
    .B(net5118),
    .Y(_04375_));
 XOR2x2_ASAP7_75t_R _10464_ (.A(net4669),
    .B(net4943),
    .Y(_04376_));
 AND2x2_ASAP7_75t_R _10465_ (.A(_04375_),
    .B(_04376_),
    .Y(_04377_));
 AND3x1_ASAP7_75t_R _10466_ (.A(net4723),
    .B(net4940),
    .C(net4939),
    .Y(_04378_));
 XOR2x2_ASAP7_75t_R _10467_ (.A(_04378_),
    .B(net4941),
    .Y(_04379_));
 INVx1_ASAP7_75t_R _10468_ (.A(_04379_),
    .Y(_04380_));
 XOR2x2_ASAP7_75t_R _10469_ (.A(net4667),
    .B(net5120),
    .Y(_04381_));
 NOR2x1_ASAP7_75t_R _10470_ (.A(net4668),
    .B(net4610),
    .Y(_04382_));
 AND2x2_ASAP7_75t_R _10471_ (.A(_04382_),
    .B(_04345_),
    .Y(_04383_));
 AND4x1_ASAP7_75t_R _10472_ (.A(net4517),
    .B(_04377_),
    .C(net4553),
    .D(_04383_),
    .Y(_04384_));
 NOR2x1_ASAP7_75t_R _10473_ (.A(net5117),
    .B(net4669),
    .Y(_04385_));
 NAND2x1_ASAP7_75t_R _10474_ (.A(net4944),
    .B(net4609),
    .Y(_04386_));
 XOR2x2_ASAP7_75t_R _10475_ (.A(_04386_),
    .B(net4945),
    .Y(_04387_));
 NOR2x1_ASAP7_75t_R _10476_ (.A(net4881),
    .B(net4612),
    .Y(_04388_));
 XOR2x2_ASAP7_75t_R _10477_ (.A(_04388_),
    .B(net5138),
    .Y(_04389_));
 NOR2x1_ASAP7_75t_R _10478_ (.A(net5141),
    .B(net5142),
    .Y(_04390_));
 AND4x1_ASAP7_75t_R _10479_ (.A(_04374_),
    .B(net4943),
    .C(net4942),
    .D(net4879),
    .Y(_04391_));
 XOR2x2_ASAP7_75t_R _10480_ (.A(_04391_),
    .B(net4946),
    .Y(_04392_));
 INVx1_ASAP7_75t_R _10481_ (.A(_04392_),
    .Y(_04393_));
 AND3x1_ASAP7_75t_R _10482_ (.A(_04385_),
    .B(net4946),
    .C(net4879),
    .Y(_04394_));
 XOR2x2_ASAP7_75t_R _10483_ (.A(net4551),
    .B(net5139),
    .Y(_04395_));
 AND2x2_ASAP7_75t_R _10484_ (.A(_04393_),
    .B(_04395_),
    .Y(_04396_));
 AND4x1_ASAP7_75t_R _10485_ (.A(_04384_),
    .B(net4514),
    .C(net4513),
    .D(net4360),
    .Y(_04397_));
 XOR2x2_ASAP7_75t_R _10486_ (.A(_04352_),
    .B(net4948),
    .Y(_04398_));
 AND3x1_ASAP7_75t_R _10487_ (.A(_04390_),
    .B(net4943),
    .C(net4942),
    .Y(_04399_));
 AND5x1_ASAP7_75t_R _10488_ (.A(net4948),
    .B(_04399_),
    .C(net5434),
    .D(net4947),
    .E(net4946),
    .Y(_04400_));
 NAND2x1_ASAP7_75t_R _10489_ (.A(_04374_),
    .B(_04400_),
    .Y(_04401_));
 XOR2x2_ASAP7_75t_R _10490_ (.A(net4511),
    .B(net4949),
    .Y(_04402_));
 AND2x2_ASAP7_75t_R _10491_ (.A(net4550),
    .B(_04402_),
    .Y(_04403_));
 AND4x1_ASAP7_75t_R _10492_ (.A(_04400_),
    .B(net4950),
    .C(net4949),
    .D(_04374_),
    .Y(_04404_));
 XOR2x2_ASAP7_75t_R _10493_ (.A(_04404_),
    .B(net4951),
    .Y(_04405_));
 AND5x1_ASAP7_75t_R _10494_ (.A(net4949),
    .B(_04394_),
    .C(net4948),
    .D(net5434),
    .E(net4947),
    .Y(_04406_));
 XOR2x2_ASAP7_75t_R _10495_ (.A(_04406_),
    .B(net4950),
    .Y(_04407_));
 NOR2x1_ASAP7_75t_R _10496_ (.A(_04405_),
    .B(_04407_),
    .Y(_04408_));
 AND3x1_ASAP7_75t_R _10497_ (.A(_04397_),
    .B(net4412),
    .C(net4411),
    .Y(_04409_));
 OR4x1_ASAP7_75t_R _10498_ (.A(net5133),
    .B(net5134),
    .C(net5135),
    .D(net5136),
    .Y(_04410_));
 NOR2x1_ASAP7_75t_R _10499_ (.A(_04410_),
    .B(_04401_),
    .Y(_04411_));
 XOR2x2_ASAP7_75t_R _10500_ (.A(_04411_),
    .B(net4953),
    .Y(_04412_));
 OR3x1_ASAP7_75t_R _10501_ (.A(_04352_),
    .B(net5137),
    .C(_04353_),
    .Y(_04413_));
 XOR2x2_ASAP7_75t_R _10502_ (.A(net4549),
    .B(net5133),
    .Y(_04414_));
 NOR2x1_ASAP7_75t_R _10503_ (.A(_04412_),
    .B(_04414_),
    .Y(_04415_));
 INVx1_ASAP7_75t_R _10504_ (.A(_04363_),
    .Y(_04416_));
 BUFx3_ASAP7_75t_R place2954 (.A(net5452),
    .Y(net2954));
 AO21x1_ASAP7_75t_R _10506_ (.A1(net4267),
    .A2(net4359),
    .B(net4320),
    .Y(_04418_));
 OR3x1_ASAP7_75t_R _10507_ (.A(_04413_),
    .B(net5131),
    .C(net5133),
    .Y(_04419_));
 XOR2x2_ASAP7_75t_R _10508_ (.A(_04419_),
    .B(net5130),
    .Y(_04420_));
 XOR2x2_ASAP7_75t_R _10509_ (.A(_04418_),
    .B(net4460),
    .Y(_04421_));
 INVx1_ASAP7_75t_R _10510_ (.A(_04421_),
    .Y(_04422_));
 AND4x1_ASAP7_75t_R _10511_ (.A(net4958),
    .B(net4957),
    .C(net4956),
    .D(net4955),
    .Y(_04423_));
 INVx1_ASAP7_75t_R _10512_ (.A(_04423_),
    .Y(_04424_));
 NOR2x1_ASAP7_75t_R _10513_ (.A(net5130),
    .B(net5131),
    .Y(_04425_));
 NAND2x1_ASAP7_75t_R _10514_ (.A(_04425_),
    .B(_04411_),
    .Y(_04426_));
 NOR2x1_ASAP7_75t_R _10515_ (.A(_04424_),
    .B(net4408),
    .Y(_04427_));
 XOR2x2_ASAP7_75t_R _10516_ (.A(_04427_),
    .B(net4959),
    .Y(_04428_));
 AND3x2_ASAP7_75t_R _10517_ (.A(_04356_),
    .B(net4958),
    .C(_04359_),
    .Y(_04429_));
 NAND3x1_ASAP7_75t_R _10518_ (.A(net4458),
    .B(net4960),
    .C(net4959),
    .Y(_04430_));
 AO21x1_ASAP7_75t_R _10519_ (.A1(_04429_),
    .A2(net4959),
    .B(net4960),
    .Y(_04431_));
 NAND2x1_ASAP7_75t_R _10520_ (.A(_04430_),
    .B(_04431_),
    .Y(_04432_));
 INVx1_ASAP7_75t_R _10521_ (.A(_04432_),
    .Y(_04433_));
 NOR2x1_ASAP7_75t_R _10522_ (.A(net4319),
    .B(net4318),
    .Y(_04434_));
 INVx1_ASAP7_75t_R _10523_ (.A(_04366_),
    .Y(_04435_));
 INVx1_ASAP7_75t_R _10524_ (.A(net4816),
    .Y(_04436_));
 AND3x1_ASAP7_75t_R _10525_ (.A(_04338_),
    .B(_04436_),
    .C(net4936),
    .Y(_04437_));
 AND3x1_ASAP7_75t_R _10526_ (.A(_04435_),
    .B(_04437_),
    .C(_04341_),
    .Y(_04438_));
 INVx1_ASAP7_75t_R _10527_ (.A(_04381_),
    .Y(_04439_));
 AND3x1_ASAP7_75t_R _10528_ (.A(_04438_),
    .B(_04380_),
    .C(_04439_),
    .Y(_04440_));
 AND2x2_ASAP7_75t_R _10529_ (.A(_04440_),
    .B(_04377_),
    .Y(_04441_));
 AND3x1_ASAP7_75t_R _10530_ (.A(_04441_),
    .B(_04372_),
    .C(_04387_),
    .Y(_04442_));
 AND2x2_ASAP7_75t_R _10531_ (.A(_04389_),
    .B(_04398_),
    .Y(_04443_));
 AND3x1_ASAP7_75t_R _10532_ (.A(_04442_),
    .B(_04396_),
    .C(_04443_),
    .Y(_04444_));
 INVx1_ASAP7_75t_R _10533_ (.A(_04407_),
    .Y(_04445_));
 AND2x2_ASAP7_75t_R _10534_ (.A(_04445_),
    .B(_04402_),
    .Y(_04446_));
 NOR2x1_ASAP7_75t_R _10535_ (.A(_04405_),
    .B(_04414_),
    .Y(_04447_));
 AND3x1_ASAP7_75t_R _10536_ (.A(_04444_),
    .B(_04446_),
    .C(_04447_),
    .Y(_04448_));
 OR3x1_ASAP7_75t_R _10537_ (.A(_04426_),
    .B(net5128),
    .C(net5129),
    .Y(_04449_));
 XOR2x2_ASAP7_75t_R _10538_ (.A(_04449_),
    .B(net5127),
    .Y(_04450_));
 AOI21x1_ASAP7_75t_R _10539_ (.A1(net4880),
    .A2(net4518),
    .B(net4958),
    .Y(_04451_));
 NOR2x2_ASAP7_75t_R _10540_ (.A(_04451_),
    .B(_04429_),
    .Y(_04452_));
 NOR2x1_ASAP7_75t_R _10541_ (.A(net4316),
    .B(net4404),
    .Y(_04453_));
 XOR2x2_ASAP7_75t_R _10542_ (.A(net4409),
    .B(net5129),
    .Y(_04454_));
 XOR2x2_ASAP7_75t_R _10543_ (.A(net4554),
    .B(net5128),
    .Y(_04455_));
 NOR2x1_ASAP7_75t_R _10544_ (.A(net4354),
    .B(net4509),
    .Y(_04456_));
 NOR2x1_ASAP7_75t_R _10545_ (.A(_04412_),
    .B(net4459),
    .Y(_04457_));
 NAND2x1_ASAP7_75t_R _10546_ (.A(_04456_),
    .B(_04457_),
    .Y(_04458_));
 INVx1_ASAP7_75t_R _10547_ (.A(_04458_),
    .Y(_04459_));
 AND3x1_ASAP7_75t_R _10548_ (.A(_04448_),
    .B(_04453_),
    .C(_04459_),
    .Y(_04460_));
 AOI21x1_ASAP7_75t_R _10549_ (.A1(_04434_),
    .A2(_04460_),
    .B(_04416_),
    .Y(_04461_));
 AND2x2_ASAP7_75t_R _10550_ (.A(net4358),
    .B(net4837),
    .Y(_04462_));
 NAND2x1_ASAP7_75t_R _10551_ (.A(net4959),
    .B(net4358),
    .Y(_04463_));
 OA21x2_ASAP7_75t_R _10552_ (.A1(_04463_),
    .A2(net5126),
    .B(net5125),
    .Y(_04464_));
 NOR2x1_ASAP7_75t_R _10553_ (.A(_04462_),
    .B(_04464_),
    .Y(_04465_));
 INVx1_ASAP7_75t_R _10554_ (.A(net4205),
    .Y(_04466_));
 XOR2x2_ASAP7_75t_R _10555_ (.A(_04461_),
    .B(_04466_),
    .Y(_04467_));
 INVx1_ASAP7_75t_R _10556_ (.A(_04467_),
    .Y(_04468_));
 NOR2x1_ASAP7_75t_R _10557_ (.A(net4318),
    .B(net4361),
    .Y(_04469_));
 AND2x2_ASAP7_75t_R _10558_ (.A(net4516),
    .B(net4553),
    .Y(_04470_));
 AND3x1_ASAP7_75t_R _10559_ (.A(net4517),
    .B(net4611),
    .C(_04470_),
    .Y(_04471_));
 AND5x1_ASAP7_75t_R _10560_ (.A(net4671),
    .B(_04471_),
    .C(net4613),
    .D(net4614),
    .E(net4552),
    .Y(_04472_));
 NOR2x1_ASAP7_75t_R _10561_ (.A(_04454_),
    .B(_04420_),
    .Y(_04473_));
 AND2x2_ASAP7_75t_R _10562_ (.A(_04473_),
    .B(_04415_),
    .Y(_04474_));
 NOR2x1_ASAP7_75t_R _10563_ (.A(_04428_),
    .B(_04452_),
    .Y(_04475_));
 NOR2x1_ASAP7_75t_R _10564_ (.A(_04455_),
    .B(_04450_),
    .Y(_04476_));
 AND2x2_ASAP7_75t_R _10565_ (.A(_04475_),
    .B(_04476_),
    .Y(_04477_));
 AND2x2_ASAP7_75t_R _10566_ (.A(net4413),
    .B(net4514),
    .Y(_04478_));
 AND3x1_ASAP7_75t_R _10567_ (.A(_04478_),
    .B(net4513),
    .C(net4512),
    .Y(_04479_));
 AND2x2_ASAP7_75t_R _10568_ (.A(_04408_),
    .B(_04403_),
    .Y(_04480_));
 AND4x1_ASAP7_75t_R _10569_ (.A(_04474_),
    .B(_04477_),
    .C(_04479_),
    .D(_04480_),
    .Y(_04481_));
 NAND2x1_ASAP7_75t_R _10570_ (.A(_04472_),
    .B(_04481_),
    .Y(_04482_));
 NOR2x1_ASAP7_75t_R _10571_ (.A(net4318),
    .B(_04482_),
    .Y(_04483_));
 AND2x2_ASAP7_75t_R _10572_ (.A(_04482_),
    .B(net4318),
    .Y(_04484_));
 OAI21x1_ASAP7_75t_R _10573_ (.A1(_04483_),
    .A2(_04484_),
    .B(net4361),
    .Y(_04485_));
 INVx1_ASAP7_75t_R _10574_ (.A(_04485_),
    .Y(_04486_));
 AOI21x1_ASAP7_75t_R _10575_ (.A1(net4837),
    .A2(net4458),
    .B(net4962),
    .Y(_04487_));
 AND3x1_ASAP7_75t_R _10576_ (.A(net4458),
    .B(net4962),
    .C(net4837),
    .Y(_04488_));
 NOR2x1_ASAP7_75t_R _10577_ (.A(_04487_),
    .B(_04488_),
    .Y(_04489_));
 NOR2x1_ASAP7_75t_R _10578_ (.A(net4205),
    .B(net4350),
    .Y(_04490_));
 NAND3x1_ASAP7_75t_R _10579_ (.A(_04460_),
    .B(_04490_),
    .C(_04434_),
    .Y(_04491_));
 NOR2x1_ASAP7_75t_R _10580_ (.A(net5127),
    .B(net4356),
    .Y(_04492_));
 AOI21x1_ASAP7_75t_R _10581_ (.A1(_04358_),
    .A2(_04492_),
    .B(net4963),
    .Y(_04493_));
 AND3x1_ASAP7_75t_R _10582_ (.A(_04492_),
    .B(net4963),
    .C(_04358_),
    .Y(_04494_));
 NOR2x1_ASAP7_75t_R _10583_ (.A(_04493_),
    .B(_04494_),
    .Y(_04495_));
 NOR2x1_ASAP7_75t_R _10584_ (.A(_04495_),
    .B(_04489_),
    .Y(_04496_));
 NOR2x1_ASAP7_75t_R _10585_ (.A(_04465_),
    .B(_04433_),
    .Y(_04497_));
 NAND3x1_ASAP7_75t_R _10586_ (.A(_04496_),
    .B(_04497_),
    .C(_04477_),
    .Y(_04498_));
 AND2x2_ASAP7_75t_R _10587_ (.A(_04479_),
    .B(net4403),
    .Y(_04499_));
 NAND2x1_ASAP7_75t_R _10588_ (.A(net4515),
    .B(_04499_),
    .Y(_04500_));
 NAND3x1_ASAP7_75t_R _10589_ (.A(net4351),
    .B(net4315),
    .C(net4359),
    .Y(_04501_));
 NOR3x1_ASAP7_75t_R _10590_ (.A(_04498_),
    .B(_04500_),
    .C(_04501_),
    .Y(_04502_));
 NAND3x1_ASAP7_75t_R _10591_ (.A(_04491_),
    .B(net4361),
    .C(_04502_),
    .Y(_04503_));
 OAI21x1_ASAP7_75t_R _10592_ (.A1(_04469_),
    .A2(_04486_),
    .B(_04503_),
    .Y(_04504_));
 NOR2x1_ASAP7_75t_R _10593_ (.A(_04468_),
    .B(_04504_),
    .Y(_04505_));
 INVx2_ASAP7_75t_R _10594_ (.A(_04505_),
    .Y(_04506_));
 INVx1_ASAP7_75t_R _10595_ (.A(net4204),
    .Y(_04507_));
 AO21x1_ASAP7_75t_R _10596_ (.A1(net4072),
    .A2(net4363),
    .B(_04507_),
    .Y(_04508_));
 NAND3x1_ASAP7_75t_R _10597_ (.A(net4072),
    .B(net4363),
    .C(_04507_),
    .Y(_04509_));
 NOR2x1_ASAP7_75t_R _10598_ (.A(net4350),
    .B(net4361),
    .Y(_04510_));
 AND3x1_ASAP7_75t_R _10599_ (.A(net4513),
    .B(net4512),
    .C(net4412),
    .Y(_04511_));
 AND3x1_ASAP7_75t_R _10600_ (.A(_04511_),
    .B(net4411),
    .C(net4359),
    .Y(_04512_));
 INVx1_ASAP7_75t_R _10601_ (.A(_04512_),
    .Y(_04513_));
 AND2x2_ASAP7_75t_R _10602_ (.A(net4315),
    .B(_04476_),
    .Y(_04514_));
 NAND3x1_ASAP7_75t_R _10603_ (.A(net4131),
    .B(_04514_),
    .C(net4264),
    .Y(_04515_));
 NOR2x1_ASAP7_75t_R _10604_ (.A(_04513_),
    .B(_04515_),
    .Y(_04516_));
 INVx1_ASAP7_75t_R _10605_ (.A(net4350),
    .Y(_04517_));
 AND5x1_ASAP7_75t_R _10606_ (.A(net4517),
    .B(net4352),
    .C(net4611),
    .D(net4552),
    .E(net4457),
    .Y(_04518_));
 AND2x2_ASAP7_75t_R _10607_ (.A(_04518_),
    .B(net4555),
    .Y(_04519_));
 AND3x1_ASAP7_75t_R _10608_ (.A(_04516_),
    .B(_04517_),
    .C(_04519_),
    .Y(_04520_));
 AOI21x1_ASAP7_75t_R _10609_ (.A1(_04519_),
    .A2(_04516_),
    .B(net4314),
    .Y(_04521_));
 OA21x2_ASAP7_75t_R _10610_ (.A1(_04520_),
    .A2(_04521_),
    .B(net4361),
    .Y(_04522_));
 AOI211x1_ASAP7_75t_R _10611_ (.A1(_04508_),
    .A2(_04509_),
    .B(_04510_),
    .C(_04522_),
    .Y(_04523_));
 NAND2x1_ASAP7_75t_R _10612_ (.A(net4361),
    .B(net4072),
    .Y(_04524_));
 AND3x1_ASAP7_75t_R _10613_ (.A(_04524_),
    .B(net4363),
    .C(net4036),
    .Y(_04525_));
 NOR2x1_ASAP7_75t_R _10614_ (.A(_04416_),
    .B(_04460_),
    .Y(_04526_));
 XNOR2x2_ASAP7_75t_R _10615_ (.A(net4319),
    .B(_04526_),
    .Y(_04527_));
 INVx1_ASAP7_75t_R _10616_ (.A(_04527_),
    .Y(_04528_));
 AOI211x1_ASAP7_75t_R _10617_ (.A1(_04506_),
    .A2(_04523_),
    .B(net4009),
    .C(net4007),
    .Y(_04529_));
 INVx1_ASAP7_75t_R _10618_ (.A(net3960),
    .Y(_04530_));
 NAND2x1_ASAP7_75t_R _10619_ (.A(_04509_),
    .B(_04508_),
    .Y(_04531_));
 NOR2x1_ASAP7_75t_R _10620_ (.A(_04510_),
    .B(_04522_),
    .Y(_04532_));
 NAND2x1_ASAP7_75t_R _10621_ (.A(_04531_),
    .B(_04532_),
    .Y(_04533_));
 NOR3x1_ASAP7_75t_R _10622_ (.A(net3988),
    .B(net4011),
    .C(_04528_),
    .Y(_04534_));
 INVx1_ASAP7_75t_R _10623_ (.A(_04525_),
    .Y(_04535_));
 OAI21x1_ASAP7_75t_R _10624_ (.A1(_04533_),
    .A2(_04534_),
    .B(_04535_),
    .Y(_04536_));
 NAND2x1_ASAP7_75t_R _10625_ (.A(net4008),
    .B(_04536_),
    .Y(_04537_));
 NAND2x1_ASAP7_75t_R _10626_ (.A(_04530_),
    .B(_04537_),
    .Y(_04538_));
 INVx1_ASAP7_75t_R _10627_ (.A(net3943),
    .Y(_04539_));
 OAI21x1_ASAP7_75t_R _10628_ (.A1(net4007),
    .A2(_04506_),
    .B(_04523_),
    .Y(_04540_));
 AOI21x1_ASAP7_75t_R _10629_ (.A1(_04535_),
    .A2(_04540_),
    .B(net4035),
    .Y(_04541_));
 INVx1_ASAP7_75t_R _10630_ (.A(net3987),
    .Y(_04542_));
 OAI21x1_ASAP7_75t_R _10631_ (.A1(_04529_),
    .A2(_04541_),
    .B(_04542_),
    .Y(_04543_));
 INVx1_ASAP7_75t_R _10632_ (.A(net3986),
    .Y(_04544_));
 INVx1_ASAP7_75t_R _10633_ (.A(net4010),
    .Y(_04545_));
 NOR2x1_ASAP7_75t_R _10634_ (.A(net4037),
    .B(_04545_),
    .Y(_04546_));
 INVx1_ASAP7_75t_R _10635_ (.A(_04546_),
    .Y(_04547_));
 NOR3x1_ASAP7_75t_R _10636_ (.A(_04536_),
    .B(_04544_),
    .C(_04547_),
    .Y(_04548_));
 AND2x2_ASAP7_75t_R _10637_ (.A(_04531_),
    .B(net4010),
    .Y(_04549_));
 AND2x2_ASAP7_75t_R _10638_ (.A(_04540_),
    .B(_04549_),
    .Y(_04550_));
 AND2x2_ASAP7_75t_R _10639_ (.A(_04409_),
    .B(net4359),
    .Y(_04551_));
 INVx1_ASAP7_75t_R _10640_ (.A(_04551_),
    .Y(_04552_));
 OR5x1_ASAP7_75t_R _10641_ (.A(net4316),
    .B(_04552_),
    .C(net4509),
    .D(net4460),
    .E(net4355),
    .Y(_04553_));
 NAND2x1_ASAP7_75t_R _10642_ (.A(net4361),
    .B(_04553_),
    .Y(_04554_));
 XOR2x2_ASAP7_75t_R _10643_ (.A(_04554_),
    .B(net4404),
    .Y(_04555_));
 INVx1_ASAP7_75t_R _10644_ (.A(_04555_),
    .Y(_04556_));
 AOI211x1_ASAP7_75t_R _10645_ (.A1(net3942),
    .A2(net3959),
    .B(net3949),
    .C(net3993),
    .Y(_04557_));
 INVx1_ASAP7_75t_R _10646_ (.A(_04550_),
    .Y(_04558_));
 OAI21x1_ASAP7_75t_R _10647_ (.A1(_04556_),
    .A2(_04543_),
    .B(_04548_),
    .Y(_04559_));
 AOI21x1_ASAP7_75t_R _10648_ (.A1(_04558_),
    .A2(net3930),
    .B(net4006),
    .Y(_04560_));
 AO21x1_ASAP7_75t_R _10649_ (.A1(net4266),
    .A2(net4206),
    .B(net4320),
    .Y(_04561_));
 XOR2x2_ASAP7_75t_R _10650_ (.A(_04561_),
    .B(net4316),
    .Y(_04562_));
 OAI21x1_ASAP7_75t_R _10651_ (.A1(_04557_),
    .A2(_04560_),
    .B(_04562_),
    .Y(_04563_));
 NOR2x1_ASAP7_75t_R _10652_ (.A(_04539_),
    .B(_04563_),
    .Y(_04564_));
 INVx1_ASAP7_75t_R _10653_ (.A(_04564_),
    .Y(_04565_));
 OAI22x1_ASAP7_75t_R _10654_ (.A1(net3942),
    .A2(net3993),
    .B1(net3959),
    .B2(net3949),
    .Y(_04566_));
 AND3x1_ASAP7_75t_R _10655_ (.A(_04536_),
    .B(net4035),
    .C(_04542_),
    .Y(_04567_));
 OAI21x1_ASAP7_75t_R _10656_ (.A1(net3977),
    .A2(_04567_),
    .B(net3994),
    .Y(_04568_));
 XOR2x2_ASAP7_75t_R _10657_ (.A(_04566_),
    .B(_04568_),
    .Y(_04569_));
 NAND2x1_ASAP7_75t_R _10658_ (.A(_04558_),
    .B(_04559_),
    .Y(_04570_));
 INVx1_ASAP7_75t_R _10659_ (.A(_04570_),
    .Y(_04571_));
 AOI21x1_ASAP7_75t_R _10660_ (.A1(_04530_),
    .A2(_04537_),
    .B(_04556_),
    .Y(_04572_));
 NOR2x1_ASAP7_75t_R _10661_ (.A(net4265),
    .B(net3995),
    .Y(_04573_));
 NOR2x1_ASAP7_75t_R _10662_ (.A(net4035),
    .B(net3987),
    .Y(_04574_));
 AOI21x1_ASAP7_75t_R _10663_ (.A1(_04573_),
    .A2(net4035),
    .B(_04574_),
    .Y(_04575_));
 INVx1_ASAP7_75t_R _10664_ (.A(_04575_),
    .Y(_04576_));
 NOR2x1_ASAP7_75t_R _10665_ (.A(net3987),
    .B(net3969),
    .Y(_04577_));
 AOI21x1_ASAP7_75t_R _10666_ (.A1(net3969),
    .A2(net3958),
    .B(_04577_),
    .Y(_04578_));
 NAND2x1_ASAP7_75t_R _10667_ (.A(_04572_),
    .B(_04578_),
    .Y(_04579_));
 NAND2x1_ASAP7_75t_R _10668_ (.A(_04576_),
    .B(net3969),
    .Y(_04580_));
 OAI21x1_ASAP7_75t_R _10669_ (.A1(net3987),
    .A2(net3969),
    .B(_04580_),
    .Y(_04581_));
 OAI21x1_ASAP7_75t_R _10670_ (.A1(net3960),
    .A2(net3950),
    .B(net4006),
    .Y(_04582_));
 NAND2x1_ASAP7_75t_R _10671_ (.A(_04581_),
    .B(_04582_),
    .Y(_04583_));
 AND2x2_ASAP7_75t_R _10672_ (.A(_04579_),
    .B(_04583_),
    .Y(_04584_));
 NAND3x1_ASAP7_75t_R _10673_ (.A(net3931),
    .B(net3941),
    .C(net3940),
    .Y(_04585_));
 OAI21x1_ASAP7_75t_R _10674_ (.A1(_04571_),
    .A2(_04584_),
    .B(_04585_),
    .Y(_04586_));
 NOR2x2_ASAP7_75t_R _10675_ (.A(net3919),
    .B(_04586_),
    .Y(_04587_));
 INVx1_ASAP7_75t_R _10676_ (.A(net3910),
    .Y(_04588_));
 AO21x1_ASAP7_75t_R _10677_ (.A1(net3900),
    .A2(net3943),
    .B(net3901),
    .Y(_04589_));
 INVx1_ASAP7_75t_R _10678_ (.A(net3931),
    .Y(_04590_));
 NAND2x1_ASAP7_75t_R _10679_ (.A(net3979),
    .B(_04572_),
    .Y(_04591_));
 AND2x2_ASAP7_75t_R _10680_ (.A(_04568_),
    .B(_04591_),
    .Y(_04592_));
 AOI21x1_ASAP7_75t_R _10681_ (.A1(net4035),
    .A2(net3981),
    .B(net3980),
    .Y(_04593_));
 NOR2x1_ASAP7_75t_R _10682_ (.A(net3978),
    .B(_04593_),
    .Y(_04594_));
 AOI21x1_ASAP7_75t_R _10683_ (.A1(_04570_),
    .A2(_04592_),
    .B(_04594_),
    .Y(_04595_));
 NOR2x1_ASAP7_75t_R _10684_ (.A(_04590_),
    .B(_04595_),
    .Y(_04596_));
 INVx1_ASAP7_75t_R _10685_ (.A(_04596_),
    .Y(_04597_));
 OA21x2_ASAP7_75t_R _10686_ (.A1(_04589_),
    .A2(_04597_),
    .B(net3919),
    .Y(_04598_));
 AOI21x1_ASAP7_75t_R _10687_ (.A1(net3886),
    .A2(net3885),
    .B(_04598_),
    .Y(_04599_));
 OAI21x1_ASAP7_75t_R _10688_ (.A1(net3899),
    .A2(_04587_),
    .B(_04565_),
    .Y(_04600_));
 AOI22x1_ASAP7_75t_R _10689_ (.A1(net3931),
    .A2(net3941),
    .B1(_04579_),
    .B2(_04583_),
    .Y(_04601_));
 NOR2x1_ASAP7_75t_R _10690_ (.A(net3948),
    .B(_04570_),
    .Y(_04602_));
 NOR2x1_ASAP7_75t_R _10691_ (.A(_04601_),
    .B(_04602_),
    .Y(_04603_));
 XOR2x2_ASAP7_75t_R _10692_ (.A(_04600_),
    .B(net3898),
    .Y(_04604_));
 XOR2x2_ASAP7_75t_R _10693_ (.A(_04538_),
    .B(net4006),
    .Y(_04605_));
 NAND2x1_ASAP7_75t_R _10694_ (.A(_04605_),
    .B(_04570_),
    .Y(_04606_));
 OAI21x1_ASAP7_75t_R _10695_ (.A1(net3933),
    .A2(net3918),
    .B(_04606_),
    .Y(_04607_));
 XOR2x2_ASAP7_75t_R _10696_ (.A(_04607_),
    .B(_04588_),
    .Y(_04608_));
 INVx1_ASAP7_75t_R _10697_ (.A(_04569_),
    .Y(_04609_));
 NAND2x1_ASAP7_75t_R _10698_ (.A(_04609_),
    .B(_04603_),
    .Y(_04610_));
 OAI21x1_ASAP7_75t_R _10699_ (.A1(_04564_),
    .A2(_04610_),
    .B(_04597_),
    .Y(_04611_));
 NAND2x1_ASAP7_75t_R _10700_ (.A(_04608_),
    .B(_04611_),
    .Y(_04612_));
 AOI21x1_ASAP7_75t_R _10701_ (.A1(_04587_),
    .A2(_04565_),
    .B(net3899),
    .Y(_04613_));
 NAND2x1_ASAP7_75t_R _10702_ (.A(net3897),
    .B(_04613_),
    .Y(_04614_));
 NAND2x1_ASAP7_75t_R _10703_ (.A(_04612_),
    .B(_04614_),
    .Y(_04615_));
 NOR2x1_ASAP7_75t_R _10704_ (.A(_04604_),
    .B(_04615_),
    .Y(_04616_));
 NOR2x1_ASAP7_75t_R _10705_ (.A(net3932),
    .B(net3920),
    .Y(_04617_));
 AOI21x1_ASAP7_75t_R _10706_ (.A1(net4071),
    .A2(_04611_),
    .B(_04617_),
    .Y(_04618_));
 AO21x1_ASAP7_75t_R _10707_ (.A1(_04551_),
    .A2(net4315),
    .B(net4320),
    .Y(_04619_));
 XOR2x2_ASAP7_75t_R _10708_ (.A(_04619_),
    .B(net4509),
    .Y(_04620_));
 INVx1_ASAP7_75t_R _10709_ (.A(net4071),
    .Y(_04621_));
 NAND2x1_ASAP7_75t_R _10710_ (.A(_04621_),
    .B(_04613_),
    .Y(_04622_));
 NAND3x1_ASAP7_75t_R _10711_ (.A(_04618_),
    .B(_04620_),
    .C(_04622_),
    .Y(_04623_));
 OAI21x1_ASAP7_75t_R _10712_ (.A1(net3868),
    .A2(net3843),
    .B(net3856),
    .Y(_04624_));
 INVx1_ASAP7_75t_R _10713_ (.A(net3897),
    .Y(_04625_));
 NOR2x1_ASAP7_75t_R _10714_ (.A(_04625_),
    .B(net3874),
    .Y(_04626_));
 XOR2x2_ASAP7_75t_R _10715_ (.A(net3897),
    .B(net3910),
    .Y(_04627_));
 NOR2x1_ASAP7_75t_R _10716_ (.A(_04627_),
    .B(net3873),
    .Y(_04628_));
 NOR2x1_ASAP7_75t_R _10717_ (.A(_04626_),
    .B(_04628_),
    .Y(_04629_));
 XOR2x2_ASAP7_75t_R _10718_ (.A(_04624_),
    .B(net3855),
    .Y(_04630_));
 XOR2x2_ASAP7_75t_R _10719_ (.A(_04617_),
    .B(_04621_),
    .Y(_04631_));
 NAND2x1_ASAP7_75t_R _10720_ (.A(_04631_),
    .B(net3874),
    .Y(_04632_));
 OAI21x1_ASAP7_75t_R _10721_ (.A1(net3909),
    .A2(net3874),
    .B(_04632_),
    .Y(_04633_));
 AOI21x1_ASAP7_75t_R _10722_ (.A1(_04623_),
    .A2(_04616_),
    .B(_04599_),
    .Y(_04634_));
 NAND2x2_ASAP7_75t_R _10723_ (.A(net3854),
    .B(_04634_),
    .Y(_04635_));
 NAND2x1_ASAP7_75t_R _10724_ (.A(net4034),
    .B(net3874),
    .Y(_04636_));
 NAND2x1_ASAP7_75t_R _10725_ (.A(net4071),
    .B(net3873),
    .Y(_04637_));
 INVx1_ASAP7_75t_R _10726_ (.A(_04620_),
    .Y(_04638_));
 AOI21x1_ASAP7_75t_R _10727_ (.A1(_04636_),
    .A2(_04637_),
    .B(_04638_),
    .Y(_04639_));
 XOR2x2_ASAP7_75t_R _10728_ (.A(_04639_),
    .B(_04633_),
    .Y(_04640_));
 XOR2x2_ASAP7_75t_R _10729_ (.A(net3875),
    .B(net3901),
    .Y(_04641_));
 NAND2x1_ASAP7_75t_R _10730_ (.A(_04641_),
    .B(_04629_),
    .Y(_04642_));
 INVx1_ASAP7_75t_R _10731_ (.A(net3909),
    .Y(_04643_));
 OAI21x1_ASAP7_75t_R _10732_ (.A1(net4034),
    .A2(net3873),
    .B(_04643_),
    .Y(_04644_));
 NOR2x1_ASAP7_75t_R _10733_ (.A(net4071),
    .B(net3874),
    .Y(_04645_));
 NOR3x1_ASAP7_75t_R _10734_ (.A(_04644_),
    .B(_04645_),
    .C(_04638_),
    .Y(_04646_));
 INVx1_ASAP7_75t_R _10735_ (.A(_04599_),
    .Y(_04647_));
 OAI21x1_ASAP7_75t_R _10736_ (.A1(_04642_),
    .A2(_04646_),
    .B(_04647_),
    .Y(_04648_));
 NAND2x1_ASAP7_75t_R _10737_ (.A(_04640_),
    .B(_04648_),
    .Y(_04649_));
 NAND2x2_ASAP7_75t_R _10738_ (.A(_04635_),
    .B(_04649_),
    .Y(_04650_));
 NOR2x2_ASAP7_75t_R _10739_ (.A(_04630_),
    .B(_04650_),
    .Y(_04651_));
 AO21x1_ASAP7_75t_R _10740_ (.A1(net3856),
    .A2(net3855),
    .B(_04641_),
    .Y(_04652_));
 NAND2x1_ASAP7_75t_R _10741_ (.A(net3856),
    .B(net3843),
    .Y(_04653_));
 NAND2x1_ASAP7_75t_R _10742_ (.A(net3867),
    .B(net3853),
    .Y(_04654_));
 OA211x2_ASAP7_75t_R _10743_ (.A1(_04652_),
    .A2(net3853),
    .B(_04653_),
    .C(_04654_),
    .Y(_04655_));
 AO21x1_ASAP7_75t_R _10744_ (.A1(net4266),
    .A2(net4353),
    .B(net4320),
    .Y(_04656_));
 XOR2x2_ASAP7_75t_R _10745_ (.A(_04656_),
    .B(net4355),
    .Y(_04657_));
 NAND2x1_ASAP7_75t_R _10746_ (.A(net4070),
    .B(_04634_),
    .Y(_04658_));
 NAND2x1_ASAP7_75t_R _10747_ (.A(net4033),
    .B(_04648_),
    .Y(_04659_));
 NAND2x1_ASAP7_75t_R _10748_ (.A(net3866),
    .B(net3865),
    .Y(_04660_));
 INVx1_ASAP7_75t_R _10749_ (.A(_04660_),
    .Y(_04661_));
 AOI21x1_ASAP7_75t_R _10750_ (.A1(_04658_),
    .A2(_04659_),
    .B(_04661_),
    .Y(_04662_));
 NAND2x1_ASAP7_75t_R _10751_ (.A(_04657_),
    .B(_04662_),
    .Y(_04663_));
 OAI21x1_ASAP7_75t_R _10752_ (.A1(_04651_),
    .A2(_04655_),
    .B(net3785),
    .Y(_04664_));
 XOR2x2_ASAP7_75t_R _10753_ (.A(_04664_),
    .B(net3802),
    .Y(_04665_));
 NOR2x1_ASAP7_75t_R _10754_ (.A(net4070),
    .B(_04634_),
    .Y(_04666_));
 NOR2x1_ASAP7_75t_R _10755_ (.A(net4033),
    .B(_04648_),
    .Y(_04667_));
 OAI21x1_ASAP7_75t_R _10756_ (.A1(net3811),
    .A2(_04667_),
    .B(_04657_),
    .Y(_04668_));
 XOR2x2_ASAP7_75t_R _10757_ (.A(_04660_),
    .B(net4033),
    .Y(_04669_));
 NAND2x1_ASAP7_75t_R _10758_ (.A(_04660_),
    .B(_04634_),
    .Y(_04670_));
 OAI21x1_ASAP7_75t_R _10759_ (.A1(net3823),
    .A2(_04669_),
    .B(_04670_),
    .Y(_04671_));
 XOR2x2_ASAP7_75t_R _10760_ (.A(_04668_),
    .B(_04671_),
    .Y(_04672_));
 AOI21x1_ASAP7_75t_R _10761_ (.A1(_04651_),
    .A2(_04663_),
    .B(_04655_),
    .Y(_04673_));
 NOR2x1_ASAP7_75t_R _10762_ (.A(_04672_),
    .B(_04673_),
    .Y(_04674_));
 INVx1_ASAP7_75t_R _10763_ (.A(net3801),
    .Y(_04675_));
 INVx1_ASAP7_75t_R _10764_ (.A(_04651_),
    .Y(_04676_));
 INVx1_ASAP7_75t_R _10765_ (.A(net4129),
    .Y(_04677_));
 OAI21x1_ASAP7_75t_R _10766_ (.A1(_04666_),
    .A2(_04667_),
    .B(net3852),
    .Y(_04678_));
 NOR2x1_ASAP7_75t_R _10767_ (.A(_04677_),
    .B(_04678_),
    .Y(_04679_));
 AO21x1_ASAP7_75t_R _10768_ (.A1(_04652_),
    .A2(_04653_),
    .B(net3824),
    .Y(_04680_));
 NAND2x1_ASAP7_75t_R _10769_ (.A(net3842),
    .B(_04680_),
    .Y(_04681_));
 OAI21x1_ASAP7_75t_R _10770_ (.A1(_04676_),
    .A2(_04679_),
    .B(_04681_),
    .Y(_04682_));
 NOR2x1_ASAP7_75t_R _10771_ (.A(_04675_),
    .B(_04682_),
    .Y(_04683_));
 NOR2x1_ASAP7_75t_R _10772_ (.A(_04674_),
    .B(_04683_),
    .Y(_04684_));
 NAND2x1_ASAP7_75t_R _10773_ (.A(_04665_),
    .B(_04684_),
    .Y(_04685_));
 AOI211x1_ASAP7_75t_R _10774_ (.A1(net3786),
    .A2(net3800),
    .B(net3813),
    .C(net4069),
    .Y(_04686_));
 NAND2x1_ASAP7_75t_R _10775_ (.A(net3786),
    .B(_04663_),
    .Y(_04687_));
 AOI21x1_ASAP7_75t_R _10776_ (.A1(_04681_),
    .A2(_04687_),
    .B(net4130),
    .Y(_04688_));
 NOR2x1_ASAP7_75t_R _10777_ (.A(net3812),
    .B(net3810),
    .Y(_04689_));
 INVx1_ASAP7_75t_R _10778_ (.A(_04689_),
    .Y(_04690_));
 OAI21x1_ASAP7_75t_R _10779_ (.A1(_04686_),
    .A2(_04688_),
    .B(_04690_),
    .Y(_04691_));
 NOR2x1_ASAP7_75t_R _10780_ (.A(_04422_),
    .B(_04691_),
    .Y(_04692_));
 AOI211x1_ASAP7_75t_R _10781_ (.A1(_04681_),
    .A2(net3814),
    .B(_04679_),
    .C(net3802),
    .Y(_04693_));
 XNOR2x2_ASAP7_75t_R _10782_ (.A(net3814),
    .B(_04693_),
    .Y(_04694_));
 INVx1_ASAP7_75t_R _10783_ (.A(_04694_),
    .Y(_04695_));
 OAI21x1_ASAP7_75t_R _10784_ (.A1(_04685_),
    .A2(_04692_),
    .B(_04695_),
    .Y(_04696_));
 NAND2x1_ASAP7_75t_R _10785_ (.A(net4073),
    .B(_04696_),
    .Y(_04697_));
 XNOR2x2_ASAP7_75t_R _10786_ (.A(net3802),
    .B(_04664_),
    .Y(_04698_));
 NAND2x1_ASAP7_75t_R _10787_ (.A(net3801),
    .B(_04673_),
    .Y(_04699_));
 OAI21x1_ASAP7_75t_R _10788_ (.A1(net3766),
    .A2(net3784),
    .B(_04699_),
    .Y(_04700_));
 NOR2x1_ASAP7_75t_R _10789_ (.A(_04698_),
    .B(_04700_),
    .Y(_04701_));
 NAND2x1_ASAP7_75t_R _10790_ (.A(net4130),
    .B(_04673_),
    .Y(_04702_));
 NAND2x1_ASAP7_75t_R _10791_ (.A(net4069),
    .B(_04682_),
    .Y(_04703_));
 AOI21x1_ASAP7_75t_R _10792_ (.A1(_04702_),
    .A2(_04703_),
    .B(net3799),
    .Y(_04704_));
 NAND2x1_ASAP7_75t_R _10793_ (.A(net4132),
    .B(_04704_),
    .Y(_04705_));
 AOI21x1_ASAP7_75t_R _10794_ (.A1(_04701_),
    .A2(_04705_),
    .B(net3758),
    .Y(_04706_));
 NAND2x1_ASAP7_75t_R _10795_ (.A(net4133),
    .B(_04706_),
    .Y(_04707_));
 NAND2x1_ASAP7_75t_R _10796_ (.A(net3700),
    .B(net3699),
    .Y(_04708_));
 INVx1_ASAP7_75t_R _10797_ (.A(_04708_),
    .Y(_04709_));
 OAI21x1_ASAP7_75t_R _10798_ (.A1(_04701_),
    .A2(net3758),
    .B(_04705_),
    .Y(_04710_));
 XOR2x2_ASAP7_75t_R _10799_ (.A(_04710_),
    .B(net3738),
    .Y(_04711_));
 XOR2x2_ASAP7_75t_R _10800_ (.A(_04689_),
    .B(net4130),
    .Y(_04712_));
 NAND2x1_ASAP7_75t_R _10801_ (.A(_04690_),
    .B(net3765),
    .Y(_04713_));
 OAI21x1_ASAP7_75t_R _10802_ (.A1(net3766),
    .A2(_04712_),
    .B(_04713_),
    .Y(_04714_));
 OAI21x1_ASAP7_75t_R _10803_ (.A1(_04686_),
    .A2(_04688_),
    .B(net4132),
    .Y(_04715_));
 XNOR2x2_ASAP7_75t_R _10804_ (.A(_04714_),
    .B(_04715_),
    .Y(_04716_));
 NAND2x1_ASAP7_75t_R _10805_ (.A(_04716_),
    .B(_04696_),
    .Y(_04717_));
 NAND2x1_ASAP7_75t_R _10806_ (.A(net3750),
    .B(_04706_),
    .Y(_04718_));
 NAND2x2_ASAP7_75t_R _10807_ (.A(_04717_),
    .B(_04718_),
    .Y(_04719_));
 NOR2x2_ASAP7_75t_R _10808_ (.A(_04711_),
    .B(_04719_),
    .Y(_04720_));
 OR2x2_ASAP7_75t_R _10809_ (.A(_04700_),
    .B(_04710_),
    .Y(_04721_));
 NOR2x1_ASAP7_75t_R _10810_ (.A(net3718),
    .B(net3737),
    .Y(_04722_));
 AOI21x1_ASAP7_75t_R _10811_ (.A1(net3757),
    .A2(_04721_),
    .B(_04722_),
    .Y(_04723_));
 AND2x2_ASAP7_75t_R _10812_ (.A(net4317),
    .B(_04446_),
    .Y(_04724_));
 AO21x1_ASAP7_75t_R _10813_ (.A1(_04724_),
    .A2(net4405),
    .B(net4320),
    .Y(_04725_));
 XOR2x2_ASAP7_75t_R _10814_ (.A(_04725_),
    .B(net4410),
    .Y(_04726_));
 INVx1_ASAP7_75t_R _10815_ (.A(_04726_),
    .Y(_04727_));
 OA21x2_ASAP7_75t_R _10816_ (.A1(_04720_),
    .A2(_04723_),
    .B(net4068),
    .Y(_04728_));
 NOR2x1_ASAP7_75t_R _10817_ (.A(net4073),
    .B(_04696_),
    .Y(_04729_));
 NOR2x1_ASAP7_75t_R _10818_ (.A(net4133),
    .B(_04706_),
    .Y(_04730_));
 NAND2x1_ASAP7_75t_R _10819_ (.A(net3756),
    .B(net3751),
    .Y(_04731_));
 OAI21x1_ASAP7_75t_R _10820_ (.A1(_04729_),
    .A2(_04730_),
    .B(net3736),
    .Y(_04732_));
 AOI211x1_ASAP7_75t_R _10821_ (.A1(net3670),
    .A2(net3686),
    .B(net3687),
    .C(net4068),
    .Y(_04733_));
 NOR2x1_ASAP7_75t_R _10822_ (.A(net4320),
    .B(net4267),
    .Y(_04734_));
 XNOR2x2_ASAP7_75t_R _10823_ (.A(net4510),
    .B(_04734_),
    .Y(_04735_));
 OAI21x1_ASAP7_75t_R _10824_ (.A1(_04728_),
    .A2(_04733_),
    .B(_04735_),
    .Y(_04736_));
 OAI21x1_ASAP7_75t_R _10825_ (.A1(net3697),
    .A2(net3696),
    .B(net4128),
    .Y(_04737_));
 INVx1_ASAP7_75t_R _10826_ (.A(_04731_),
    .Y(_04738_));
 NOR2x1_ASAP7_75t_R _10827_ (.A(net4133),
    .B(_04738_),
    .Y(_04739_));
 NOR2x1_ASAP7_75t_R _10828_ (.A(net4073),
    .B(net3736),
    .Y(_04740_));
 OAI21x1_ASAP7_75t_R _10829_ (.A1(_04739_),
    .A2(_04740_),
    .B(net3709),
    .Y(_04741_));
 OAI21x1_ASAP7_75t_R _10830_ (.A1(net3717),
    .A2(net3709),
    .B(_04741_),
    .Y(_04742_));
 INVx1_ASAP7_75t_R _10831_ (.A(net3684),
    .Y(_04743_));
 AOI211x1_ASAP7_75t_R _10832_ (.A1(net3669),
    .A2(net3685),
    .B(_04743_),
    .C(net3687),
    .Y(_04744_));
 XOR2x2_ASAP7_75t_R _10833_ (.A(_04737_),
    .B(_04742_),
    .Y(_04745_));
 AOI21x1_ASAP7_75t_R _10834_ (.A1(_04697_),
    .A2(_04707_),
    .B(_04738_),
    .Y(_04746_));
 NAND2x1_ASAP7_75t_R _10835_ (.A(_04726_),
    .B(_04746_),
    .Y(_04747_));
 AOI21x1_ASAP7_75t_R _10836_ (.A1(_04720_),
    .A2(_04747_),
    .B(_04723_),
    .Y(_04748_));
 NOR2x1_ASAP7_75t_R _10837_ (.A(_04745_),
    .B(net3655),
    .Y(_04749_));
 NOR2x1_ASAP7_75t_R _10838_ (.A(_04744_),
    .B(_04749_),
    .Y(_04750_));
 OAI21x1_ASAP7_75t_R _10839_ (.A1(net3671),
    .A2(net3647),
    .B(_04750_),
    .Y(_04751_));
 INVx1_ASAP7_75t_R _10840_ (.A(_04720_),
    .Y(_04752_));
 NOR2x1_ASAP7_75t_R _10841_ (.A(_04727_),
    .B(_04732_),
    .Y(_04753_));
 INVx1_ASAP7_75t_R _10842_ (.A(_04723_),
    .Y(_04754_));
 OAI21x1_ASAP7_75t_R _10843_ (.A1(_04752_),
    .A2(_04753_),
    .B(_04754_),
    .Y(_04755_));
 INVx1_ASAP7_75t_R _10844_ (.A(_04719_),
    .Y(_04756_));
 OAI21x1_ASAP7_75t_R _10845_ (.A1(_04727_),
    .A2(_04732_),
    .B(_04756_),
    .Y(_04757_));
 NAND3x1_ASAP7_75t_R _10846_ (.A(net3683),
    .B(net4128),
    .C(net3688),
    .Y(_04758_));
 NAND2x1_ASAP7_75t_R _10847_ (.A(_04757_),
    .B(_04758_),
    .Y(_04759_));
 NOR2x1_ASAP7_75t_R _10848_ (.A(net3666),
    .B(net3687),
    .Y(_04760_));
 AOI21x1_ASAP7_75t_R _10849_ (.A1(_04755_),
    .A2(_04759_),
    .B(_04760_),
    .Y(_04761_));
 INVx1_ASAP7_75t_R _10850_ (.A(_04761_),
    .Y(_04762_));
 NAND2x1_ASAP7_75t_R _10851_ (.A(net3684),
    .B(_04748_),
    .Y(_04763_));
 OAI21x1_ASAP7_75t_R _10852_ (.A1(net3654),
    .A2(_04745_),
    .B(_04763_),
    .Y(_04764_));
 NOR2x1_ASAP7_75t_R _10853_ (.A(_04762_),
    .B(_04764_),
    .Y(_04765_));
 INVx1_ASAP7_75t_R _10854_ (.A(_04728_),
    .Y(_04766_));
 NAND2x1_ASAP7_75t_R _10855_ (.A(net4127),
    .B(_04748_),
    .Y(_04767_));
 INVx1_ASAP7_75t_R _10856_ (.A(_04735_),
    .Y(_04768_));
 AOI21x1_ASAP7_75t_R _10857_ (.A1(_04766_),
    .A2(_04767_),
    .B(_04768_),
    .Y(_04769_));
 NAND2x1_ASAP7_75t_R _10858_ (.A(net3689),
    .B(_04769_),
    .Y(_04770_));
 OAI21x1_ASAP7_75t_R _10859_ (.A1(net3667),
    .A2(_04757_),
    .B(net3698),
    .Y(_04771_));
 OAI21x1_ASAP7_75t_R _10860_ (.A1(net3698),
    .A2(net3653),
    .B(_04771_),
    .Y(_04772_));
 INVx1_ASAP7_75t_R _10861_ (.A(_04772_),
    .Y(_04773_));
 AOI21x1_ASAP7_75t_R _10862_ (.A1(_04765_),
    .A2(_04770_),
    .B(_04773_),
    .Y(_04774_));
 NOR2x1_ASAP7_75t_R _10863_ (.A(_04709_),
    .B(_04736_),
    .Y(_04775_));
 OAI21x1_ASAP7_75t_R _10864_ (.A1(net3627),
    .A2(net3626),
    .B(net3629),
    .Y(_04776_));
 OAI21x1_ASAP7_75t_R _10865_ (.A1(_04751_),
    .A2(_04774_),
    .B(_04776_),
    .Y(_04777_));
 NAND2x1_ASAP7_75t_R _10866_ (.A(net3627),
    .B(net3630),
    .Y(_04778_));
 AOI21x1_ASAP7_75t_R _10867_ (.A1(net3627),
    .A2(_04778_),
    .B(_04751_),
    .Y(_04779_));
 INVx1_ASAP7_75t_R _10868_ (.A(net3685),
    .Y(_04780_));
 AOI21x1_ASAP7_75t_R _10869_ (.A1(_04780_),
    .A2(net3645),
    .B(net3684),
    .Y(_04781_));
 NOR2x1_ASAP7_75t_R _10870_ (.A(net3668),
    .B(_04748_),
    .Y(_04782_));
 OAI21x1_ASAP7_75t_R _10871_ (.A1(_04781_),
    .A2(_04782_),
    .B(_04761_),
    .Y(_04783_));
 NOR2x1_ASAP7_75t_R _10872_ (.A(net3604),
    .B(net3626),
    .Y(_04784_));
 INVx1_ASAP7_75t_R _10873_ (.A(_04784_),
    .Y(_04785_));
 OA21x2_ASAP7_75t_R _10874_ (.A1(_04779_),
    .A2(net3630),
    .B(_04785_),
    .Y(_04786_));
 BUFx3_ASAP7_75t_R place2953 (.A(_02251_),
    .Y(net2953));
 NOR2x1_ASAP7_75t_R _10876_ (.A(net3630),
    .B(net3574),
    .Y(_04788_));
 NOR2x1_ASAP7_75t_R _10877_ (.A(net4320),
    .B(net4263),
    .Y(_04789_));
 XNOR2x2_ASAP7_75t_R _10878_ (.A(net4461),
    .B(_04789_),
    .Y(_04790_));
 OAI21x1_ASAP7_75t_R _10879_ (.A1(_04783_),
    .A2(_04775_),
    .B(_04772_),
    .Y(_04791_));
 NAND2x2_ASAP7_75t_R _10880_ (.A(net4067),
    .B(_04791_),
    .Y(_04792_));
 NAND2x1_ASAP7_75t_R _10881_ (.A(net4126),
    .B(_04774_),
    .Y(_04793_));
 NOR2x1_ASAP7_75t_R _10882_ (.A(net3657),
    .B(net3656),
    .Y(_04794_));
 AOI21x1_ASAP7_75t_R _10883_ (.A1(_04792_),
    .A2(_04793_),
    .B(_04794_),
    .Y(_04795_));
 XOR2x2_ASAP7_75t_R _10884_ (.A(_04708_),
    .B(net4127),
    .Y(_04796_));
 NOR2x1_ASAP7_75t_R _10885_ (.A(_04709_),
    .B(net3645),
    .Y(_04797_));
 AOI21x1_ASAP7_75t_R _10886_ (.A1(net3646),
    .A2(_04796_),
    .B(_04797_),
    .Y(_04798_));
 XOR2x2_ASAP7_75t_R _10887_ (.A(_04798_),
    .B(net3647),
    .Y(_04799_));
 NAND2x1_ASAP7_75t_R _10888_ (.A(_04791_),
    .B(_04799_),
    .Y(_04800_));
 INVx1_ASAP7_75t_R _10889_ (.A(net3603),
    .Y(_04801_));
 NAND2x1_ASAP7_75t_R _10890_ (.A(_04801_),
    .B(net3591),
    .Y(_04802_));
 NAND2x1_ASAP7_75t_R _10891_ (.A(_04800_),
    .B(_04802_),
    .Y(_04803_));
 AOI21x1_ASAP7_75t_R _10892_ (.A1(net4124),
    .A2(net3559),
    .B(_04803_),
    .Y(_04804_));
 OAI21x1_ASAP7_75t_R _10893_ (.A1(_04786_),
    .A2(_04788_),
    .B(_04804_),
    .Y(_04805_));
 AOI21x1_ASAP7_75t_R _10894_ (.A1(net3605),
    .A2(net3606),
    .B(net3631),
    .Y(_04806_));
 NOR2x1_ASAP7_75t_R _10895_ (.A(_04806_),
    .B(net3598),
    .Y(_04807_));
 NAND3x1_ASAP7_75t_R _10896_ (.A(_04807_),
    .B(net3571),
    .C(net3589),
    .Y(_04808_));
 AOI21x1_ASAP7_75t_R _10897_ (.A1(net4124),
    .A2(net3559),
    .B(_04808_),
    .Y(_04809_));
 AOI21x1_ASAP7_75t_R _10898_ (.A1(net3574),
    .A2(net3534),
    .B(_04809_),
    .Y(_04810_));
 INVx1_ASAP7_75t_R _10899_ (.A(_04810_),
    .Y(_04811_));
 INVx1_ASAP7_75t_R _10900_ (.A(_04786_),
    .Y(_04812_));
 NAND2x1_ASAP7_75t_R _10901_ (.A(net4124),
    .B(_04795_),
    .Y(_04813_));
 INVx1_ASAP7_75t_R _10902_ (.A(_04813_),
    .Y(_04814_));
 OAI21x1_ASAP7_75t_R _10903_ (.A1(_04812_),
    .A2(_04814_),
    .B(_04803_),
    .Y(_04815_));
 NAND2x1_ASAP7_75t_R _10904_ (.A(_04805_),
    .B(_04815_),
    .Y(_04816_));
 INVx1_ASAP7_75t_R _10905_ (.A(_04816_),
    .Y(_04817_));
 NOR2x1_ASAP7_75t_R _10906_ (.A(net3647),
    .B(_04774_),
    .Y(_04818_));
 INVx1_ASAP7_75t_R _10907_ (.A(_04818_),
    .Y(_04819_));
 INVx1_ASAP7_75t_R _10908_ (.A(_04794_),
    .Y(_04820_));
 AO21x1_ASAP7_75t_R _10909_ (.A1(_04791_),
    .A2(net4126),
    .B(_04820_),
    .Y(_04821_));
 NAND2x1_ASAP7_75t_R _10910_ (.A(_04819_),
    .B(_04821_),
    .Y(_04822_));
 INVx1_ASAP7_75t_R _10911_ (.A(_04790_),
    .Y(_04823_));
 AOI21x1_ASAP7_75t_R _10912_ (.A1(net3590),
    .A2(net3572),
    .B(_04823_),
    .Y(_04824_));
 XOR2x2_ASAP7_75t_R _10913_ (.A(_04822_),
    .B(_04824_),
    .Y(_04825_));
 OAI21x1_ASAP7_75t_R _10914_ (.A1(net3647),
    .A2(net3591),
    .B(net3603),
    .Y(_04826_));
 NAND3x1_ASAP7_75t_R _10915_ (.A(_04791_),
    .B(net3689),
    .C(net3628),
    .Y(_04827_));
 AOI21x1_ASAP7_75t_R _10916_ (.A1(_04826_),
    .A2(_04827_),
    .B(_04777_),
    .Y(_04828_));
 AOI21x1_ASAP7_75t_R _10917_ (.A1(_04828_),
    .A2(_04813_),
    .B(_04786_),
    .Y(_04829_));
 NOR2x1_ASAP7_75t_R _10918_ (.A(_04825_),
    .B(_04829_),
    .Y(_04830_));
 AOI211x1_ASAP7_75t_R _10919_ (.A1(_04813_),
    .A2(_04828_),
    .B(net3547),
    .C(_04786_),
    .Y(_04831_));
 NOR2x1_ASAP7_75t_R _10920_ (.A(_04830_),
    .B(_04831_),
    .Y(_04832_));
 NAND2x1_ASAP7_75t_R _10921_ (.A(_04817_),
    .B(_04832_),
    .Y(_04833_));
 AOI21x1_ASAP7_75t_R _10922_ (.A1(net4321),
    .A2(net4412),
    .B(net4320),
    .Y(_04834_));
 XOR2x2_ASAP7_75t_R _10923_ (.A(_04834_),
    .B(net4406),
    .Y(_04835_));
 INVx1_ASAP7_75t_R _10924_ (.A(_04835_),
    .Y(_04836_));
 NOR2x1_ASAP7_75t_R _10925_ (.A(net4067),
    .B(_04791_),
    .Y(_04837_));
 INVx1_ASAP7_75t_R _10926_ (.A(net3590),
    .Y(_04838_));
 OAI21x1_ASAP7_75t_R _10927_ (.A1(_04837_),
    .A2(_04838_),
    .B(net3625),
    .Y(_04839_));
 AOI211x1_ASAP7_75t_R _10928_ (.A1(_04828_),
    .A2(_04839_),
    .B(_04786_),
    .C(net4066),
    .Y(_04840_));
 OAI21x1_ASAP7_75t_R _10929_ (.A1(net4066),
    .A2(_04839_),
    .B(_04828_),
    .Y(_04841_));
 AOI21x1_ASAP7_75t_R _10930_ (.A1(_04812_),
    .A2(_04841_),
    .B(net4125),
    .Y(_04842_));
 NAND2x1_ASAP7_75t_R _10931_ (.A(net3590),
    .B(net3572),
    .Y(_04843_));
 OAI21x1_ASAP7_75t_R _10932_ (.A1(_04840_),
    .A2(_04842_),
    .B(net3558),
    .Y(_04844_));
 NOR2x1_ASAP7_75t_R _10933_ (.A(_04836_),
    .B(_04844_),
    .Y(_04845_));
 AOI21x1_ASAP7_75t_R _10934_ (.A1(_04811_),
    .A2(_04833_),
    .B(net3497),
    .Y(_04846_));
 INVx1_ASAP7_75t_R _10935_ (.A(net3498),
    .Y(_04847_));
 XOR2x2_ASAP7_75t_R _10936_ (.A(_04846_),
    .B(_04847_),
    .Y(_04848_));
 XOR2x2_ASAP7_75t_R _10937_ (.A(_04843_),
    .B(net4066),
    .Y(_04849_));
 NOR2x1_ASAP7_75t_R _10938_ (.A(_04849_),
    .B(net3533),
    .Y(_04850_));
 AOI21x1_ASAP7_75t_R _10939_ (.A1(net3558),
    .A2(net3533),
    .B(_04850_),
    .Y(_04851_));
 OAI21x1_ASAP7_75t_R _10940_ (.A1(net3546),
    .A2(net3531),
    .B(net4203),
    .Y(_04852_));
 XOR2x2_ASAP7_75t_R _10941_ (.A(_04851_),
    .B(_04852_),
    .Y(_04853_));
 OAI21x1_ASAP7_75t_R _10942_ (.A1(_04845_),
    .A2(_04833_),
    .B(_04811_),
    .Y(_04854_));
 NAND2x1_ASAP7_75t_R _10943_ (.A(_04853_),
    .B(_04854_),
    .Y(_04855_));
 INVx1_ASAP7_75t_R _10944_ (.A(net3496),
    .Y(_04856_));
 NOR3x1_ASAP7_75t_R _10945_ (.A(_04816_),
    .B(net3532),
    .C(net3515),
    .Y(_04857_));
 INVx1_ASAP7_75t_R _10946_ (.A(_04840_),
    .Y(_04858_));
 OAI21x1_ASAP7_75t_R _10947_ (.A1(net3573),
    .A2(_04809_),
    .B(net4066),
    .Y(_04859_));
 INVx1_ASAP7_75t_R _10948_ (.A(net3558),
    .Y(_04860_));
 AOI21x1_ASAP7_75t_R _10949_ (.A1(_04858_),
    .A2(_04859_),
    .B(_04860_),
    .Y(_04861_));
 NAND2x1_ASAP7_75t_R _10950_ (.A(net4203),
    .B(_04861_),
    .Y(_04862_));
 AOI21x1_ASAP7_75t_R _10951_ (.A1(_04857_),
    .A2(_04862_),
    .B(net3516),
    .Y(_04863_));
 NAND2x1_ASAP7_75t_R _10952_ (.A(_04856_),
    .B(_04863_),
    .Y(_04864_));
 NAND2x2_ASAP7_75t_R _10953_ (.A(_04855_),
    .B(_04864_),
    .Y(_04865_));
 NOR2x2_ASAP7_75t_R _10954_ (.A(_04848_),
    .B(_04865_),
    .Y(_04866_));
 NOR2x1_ASAP7_75t_R _10955_ (.A(net4317),
    .B(net4320),
    .Y(_04867_));
 XOR2x2_ASAP7_75t_R _10956_ (.A(_04867_),
    .B(net4462),
    .Y(_04868_));
 NAND2x1_ASAP7_75t_R _10957_ (.A(net4123),
    .B(_04854_),
    .Y(_04869_));
 NAND2x1_ASAP7_75t_R _10958_ (.A(net4203),
    .B(_04863_),
    .Y(_04870_));
 NAND2x1_ASAP7_75t_R _10959_ (.A(net3530),
    .B(net3529),
    .Y(_04871_));
 INVx1_ASAP7_75t_R _10960_ (.A(_04871_),
    .Y(_04872_));
 AOI21x1_ASAP7_75t_R _10961_ (.A1(_04869_),
    .A2(_04870_),
    .B(_04872_),
    .Y(_04873_));
 NAND2x1_ASAP7_75t_R _10962_ (.A(_04868_),
    .B(_04873_),
    .Y(_04874_));
 NOR2x1_ASAP7_75t_R _10963_ (.A(_04847_),
    .B(net3497),
    .Y(_04875_));
 AO21x1_ASAP7_75t_R _10964_ (.A1(_04875_),
    .A2(net3516),
    .B(_04817_),
    .Y(_04876_));
 NAND2x1_ASAP7_75t_R _10965_ (.A(net3489),
    .B(net3495),
    .Y(_04877_));
 AND2x2_ASAP7_75t_R _10966_ (.A(_04876_),
    .B(_04877_),
    .Y(_04878_));
 AOI21x1_ASAP7_75t_R _10967_ (.A1(_04866_),
    .A2(_04874_),
    .B(_04878_),
    .Y(_04879_));
 NOR2x1_ASAP7_75t_R _10968_ (.A(net4123),
    .B(net3470),
    .Y(_04880_));
 NOR2x1_ASAP7_75t_R _10969_ (.A(net4202),
    .B(net3480),
    .Y(_04881_));
 OAI21x1_ASAP7_75t_R _10970_ (.A1(_04880_),
    .A2(_04881_),
    .B(_04868_),
    .Y(_04882_));
 XOR2x2_ASAP7_75t_R _10971_ (.A(_04871_),
    .B(net4202),
    .Y(_04883_));
 NAND2x1_ASAP7_75t_R _10972_ (.A(_04883_),
    .B(net3470),
    .Y(_04884_));
 OAI21x1_ASAP7_75t_R _10973_ (.A1(net3494),
    .A2(net3470),
    .B(_04884_),
    .Y(_04885_));
 XOR2x2_ASAP7_75t_R _10974_ (.A(_04882_),
    .B(_04885_),
    .Y(_04886_));
 NAND2x1_ASAP7_75t_R _10975_ (.A(net3438),
    .B(_04879_),
    .Y(_04887_));
 OAI21x1_ASAP7_75t_R _10976_ (.A1(_04879_),
    .A2(_04886_),
    .B(_04887_),
    .Y(_04888_));
 OAI21x1_ASAP7_75t_R _10977_ (.A1(_04866_),
    .A2(_04878_),
    .B(_04874_),
    .Y(_04889_));
 XOR2x2_ASAP7_75t_R _10978_ (.A(_04889_),
    .B(net3440),
    .Y(_04890_));
 INVx1_ASAP7_75t_R _10979_ (.A(_04890_),
    .Y(_04891_));
 NOR2x1_ASAP7_75t_R _10980_ (.A(_04888_),
    .B(_04891_),
    .Y(_04892_));
 NAND2x1_ASAP7_75t_R _10981_ (.A(net3455),
    .B(net3469),
    .Y(_04893_));
 NAND2x1_ASAP7_75t_R _10982_ (.A(net4201),
    .B(_04879_),
    .Y(_04894_));
 INVx1_ASAP7_75t_R _10983_ (.A(_04868_),
    .Y(_04895_));
 INVx1_ASAP7_75t_R _10984_ (.A(_04848_),
    .Y(_04896_));
 INVx1_ASAP7_75t_R _10985_ (.A(net3439),
    .Y(_04897_));
 NAND2x1_ASAP7_75t_R _10986_ (.A(_04896_),
    .B(_04897_),
    .Y(_04898_));
 OAI21x1_ASAP7_75t_R _10987_ (.A1(_04880_),
    .A2(_04881_),
    .B(net3514),
    .Y(_04899_));
 NOR2x1_ASAP7_75t_R _10988_ (.A(_04895_),
    .B(_04899_),
    .Y(_04900_));
 INVx1_ASAP7_75t_R _10989_ (.A(_04878_),
    .Y(_04901_));
 OAI21x1_ASAP7_75t_R _10990_ (.A1(_04898_),
    .A2(_04900_),
    .B(_04901_),
    .Y(_04902_));
 NAND2x1_ASAP7_75t_R _10991_ (.A(net4121),
    .B(_04902_),
    .Y(_04903_));
 OR3x1_ASAP7_75t_R _10992_ (.A(net4321),
    .B(net4416),
    .C(net4415),
    .Y(_04904_));
 XNOR2x2_ASAP7_75t_R _10993_ (.A(net4550),
    .B(_04904_),
    .Y(_04905_));
 INVx1_ASAP7_75t_R _10994_ (.A(_04905_),
    .Y(_04906_));
 AOI21x1_ASAP7_75t_R _10995_ (.A1(_04894_),
    .A2(_04903_),
    .B(_04906_),
    .Y(_04907_));
 NAND2x1_ASAP7_75t_R _10996_ (.A(net3437),
    .B(_04907_),
    .Y(_04908_));
 NAND2x1_ASAP7_75t_R _10997_ (.A(_04892_),
    .B(_04908_),
    .Y(_04909_));
 NOR2x1_ASAP7_75t_R _10998_ (.A(net3440),
    .B(_04889_),
    .Y(_04910_));
 XOR2x2_ASAP7_75t_R _10999_ (.A(_04910_),
    .B(net3436),
    .Y(_04911_));
 INVx2_ASAP7_75t_R _11000_ (.A(_04911_),
    .Y(_04912_));
 INVx1_ASAP7_75t_R _11001_ (.A(_04893_),
    .Y(_04913_));
 AOI211x1_ASAP7_75t_R _11002_ (.A1(net3422),
    .A2(_04899_),
    .B(net3454),
    .C(net4122),
    .Y(_04914_));
 OAI21x1_ASAP7_75t_R _11003_ (.A1(_04895_),
    .A2(net3435),
    .B(net3422),
    .Y(_04915_));
 AOI21x1_ASAP7_75t_R _11004_ (.A1(_04901_),
    .A2(_04915_),
    .B(net4201),
    .Y(_04916_));
 OAI21x1_ASAP7_75t_R _11005_ (.A1(_04914_),
    .A2(_04916_),
    .B(_04905_),
    .Y(_04917_));
 NOR2x2_ASAP7_75t_R _11006_ (.A(_04886_),
    .B(_04879_),
    .Y(_04918_));
 INVx1_ASAP7_75t_R _11007_ (.A(net3438),
    .Y(_04919_));
 NOR2x1_ASAP7_75t_R _11008_ (.A(_04919_),
    .B(_04902_),
    .Y(_04920_));
 NOR2x2_ASAP7_75t_R _11009_ (.A(_04918_),
    .B(_04920_),
    .Y(_04921_));
 OAI21x1_ASAP7_75t_R _11010_ (.A1(net3421),
    .A2(net3382),
    .B(net3372),
    .Y(_04922_));
 OAI21x1_ASAP7_75t_R _11011_ (.A1(_04912_),
    .A2(_04922_),
    .B(net3385),
    .Y(_04923_));
 NAND2x1_ASAP7_75t_R _11012_ (.A(_04909_),
    .B(_04923_),
    .Y(_04924_));
 INVx3_ASAP7_75t_R _11013_ (.A(_04924_),
    .Y(_04925_));
 AOI21x1_ASAP7_75t_R _11014_ (.A1(_04892_),
    .A2(_04908_),
    .B(net3383),
    .Y(_04926_));
 NOR2x1_ASAP7_75t_R _11015_ (.A(_04913_),
    .B(_04917_),
    .Y(_04927_));
 XOR2x2_ASAP7_75t_R _11016_ (.A(net3371),
    .B(net3386),
    .Y(_04928_));
 NOR2x1_ASAP7_75t_R _11017_ (.A(net3372),
    .B(net3383),
    .Y(_04929_));
 INVx1_ASAP7_75t_R _11018_ (.A(_04929_),
    .Y(_04930_));
 OAI21x1_ASAP7_75t_R _11019_ (.A1(_04926_),
    .A2(_04928_),
    .B(_04930_),
    .Y(_04931_));
 XOR2x2_ASAP7_75t_R _11020_ (.A(_04893_),
    .B(net4121),
    .Y(_04932_));
 NAND2x1_ASAP7_75t_R _11021_ (.A(_04893_),
    .B(net3410),
    .Y(_04933_));
 OAI21x1_ASAP7_75t_R _11022_ (.A1(net3410),
    .A2(_04932_),
    .B(_04933_),
    .Y(_04934_));
 XOR2x2_ASAP7_75t_R _11023_ (.A(net3382),
    .B(_04934_),
    .Y(_04935_));
 INVx1_ASAP7_75t_R _11024_ (.A(_04935_),
    .Y(_04936_));
 NAND2x1_ASAP7_75t_R _11025_ (.A(_04890_),
    .B(_04921_),
    .Y(_04937_));
 OAI21x1_ASAP7_75t_R _11026_ (.A1(_04937_),
    .A2(_04927_),
    .B(_04912_),
    .Y(_04938_));
 NAND2x1_ASAP7_75t_R _11027_ (.A(_04936_),
    .B(net3342),
    .Y(_04939_));
 NAND2x1_ASAP7_75t_R _11028_ (.A(net3381),
    .B(_04926_),
    .Y(_04940_));
 NAND2x1_ASAP7_75t_R _11029_ (.A(_04939_),
    .B(_04940_),
    .Y(_04941_));
 NOR2x1_ASAP7_75t_R _11030_ (.A(_04931_),
    .B(_04941_),
    .Y(_04942_));
 AO21x1_ASAP7_75t_R _11031_ (.A1(net4360),
    .A2(net4357),
    .B(net4320),
    .Y(_04943_));
 XNOR2x2_ASAP7_75t_R _11032_ (.A(net4513),
    .B(_04943_),
    .Y(_04944_));
 INVx1_ASAP7_75t_R _11033_ (.A(_04944_),
    .Y(_04945_));
 OAI21x1_ASAP7_75t_R _11034_ (.A1(net3311),
    .A2(_04942_),
    .B(net4119),
    .Y(_04946_));
 XOR2x2_ASAP7_75t_R _11035_ (.A(net3371),
    .B(net3372),
    .Y(_04947_));
 AOI21x1_ASAP7_75t_R _11036_ (.A1(net3343),
    .A2(_04947_),
    .B(_04929_),
    .Y(_04948_));
 NAND2x1_ASAP7_75t_R _11037_ (.A(_04935_),
    .B(net3342),
    .Y(_04949_));
 INVx1_ASAP7_75t_R _11038_ (.A(net3381),
    .Y(_04950_));
 NAND2x1_ASAP7_75t_R _11039_ (.A(_04950_),
    .B(_04926_),
    .Y(_04951_));
 NAND2x1_ASAP7_75t_R _11040_ (.A(_04949_),
    .B(_04951_),
    .Y(_04952_));
 AOI21x1_ASAP7_75t_R _11041_ (.A1(_04948_),
    .A2(_04952_),
    .B(_04925_),
    .Y(_04953_));
 NOR2x1_ASAP7_75t_R _11042_ (.A(net4120),
    .B(net3343),
    .Y(_04954_));
 AOI21x1_ASAP7_75t_R _11043_ (.A1(net3373),
    .A2(net3344),
    .B(net4200),
    .Y(_04955_));
 OAI21x1_ASAP7_75t_R _11044_ (.A1(_04954_),
    .A2(_04955_),
    .B(_04944_),
    .Y(_04956_));
 NAND2x1_ASAP7_75t_R _11045_ (.A(_04894_),
    .B(net3384),
    .Y(_04957_));
 INVx1_ASAP7_75t_R _11046_ (.A(_04957_),
    .Y(_04958_));
 NOR2x2_ASAP7_75t_R _11047_ (.A(_04958_),
    .B(net3343),
    .Y(_04959_));
 XOR2x2_ASAP7_75t_R _11048_ (.A(_04957_),
    .B(net4120),
    .Y(_04960_));
 AOI21x1_ASAP7_75t_R _11049_ (.A1(net3373),
    .A2(net3344),
    .B(_04960_),
    .Y(_04961_));
 OAI21x1_ASAP7_75t_R _11050_ (.A1(_04959_),
    .A2(_04961_),
    .B(_04924_),
    .Y(_04962_));
 NOR2x2_ASAP7_75t_R _11051_ (.A(_04956_),
    .B(_04962_),
    .Y(_04963_));
 OAI21x1_ASAP7_75t_R _11052_ (.A1(_04953_),
    .A2(_04963_),
    .B(net4199),
    .Y(_04964_));
 NAND2x1_ASAP7_75t_R _11053_ (.A(net3273),
    .B(net3272),
    .Y(_04965_));
 NOR2x1_ASAP7_75t_R _11054_ (.A(net3360),
    .B(net3308),
    .Y(_04966_));
 OAI21x1_ASAP7_75t_R _11055_ (.A1(net3328),
    .A2(_04966_),
    .B(net3310),
    .Y(_04967_));
 NOR2x1_ASAP7_75t_R _11056_ (.A(net3311),
    .B(_04931_),
    .Y(_04968_));
 NAND2x1_ASAP7_75t_R _11057_ (.A(net4120),
    .B(net3343),
    .Y(_04969_));
 NAND2x1_ASAP7_75t_R _11058_ (.A(net4200),
    .B(_04926_),
    .Y(_04970_));
 AOI21x1_ASAP7_75t_R _11059_ (.A1(_04969_),
    .A2(_04970_),
    .B(_04945_),
    .Y(_04971_));
 AOI21x1_ASAP7_75t_R _11060_ (.A1(net3370),
    .A2(_04971_),
    .B(_04941_),
    .Y(_04972_));
 OAI21x1_ASAP7_75t_R _11061_ (.A1(net3311),
    .A2(_04968_),
    .B(_04972_),
    .Y(_04973_));
 NAND2x1_ASAP7_75t_R _11062_ (.A(_04967_),
    .B(_04973_),
    .Y(_04974_));
 OAI21x1_ASAP7_75t_R _11063_ (.A1(_04931_),
    .A2(_04941_),
    .B(net3328),
    .Y(_04975_));
 OAI21x1_ASAP7_75t_R _11064_ (.A1(net3308),
    .A2(net3307),
    .B(_04975_),
    .Y(_04976_));
 NOR2x1_ASAP7_75t_R _11065_ (.A(_04959_),
    .B(_04961_),
    .Y(_04977_));
 XOR2x2_ASAP7_75t_R _11066_ (.A(_04971_),
    .B(_04977_),
    .Y(_04978_));
 INVx1_ASAP7_75t_R _11067_ (.A(net3305),
    .Y(_04979_));
 OAI21x1_ASAP7_75t_R _11068_ (.A1(_04953_),
    .A2(net3288),
    .B(_04979_),
    .Y(_04980_));
 OAI21x1_ASAP7_75t_R _11069_ (.A1(_04976_),
    .A2(_04978_),
    .B(_04980_),
    .Y(_04981_));
 NOR2x1_ASAP7_75t_R _11070_ (.A(_04974_),
    .B(_04981_),
    .Y(_04982_));
 NAND2x1_ASAP7_75t_R _11071_ (.A(net3325),
    .B(net3324),
    .Y(_04983_));
 AND2x2_ASAP7_75t_R _11072_ (.A(net4414),
    .B(net4514),
    .Y(_04984_));
 AO21x1_ASAP7_75t_R _11073_ (.A1(_04984_),
    .A2(net4413),
    .B(net4320),
    .Y(_04985_));
 XNOR2x2_ASAP7_75t_R _11074_ (.A(net4512),
    .B(_04985_),
    .Y(_04986_));
 INVx1_ASAP7_75t_R _11075_ (.A(_04986_),
    .Y(_04987_));
 AOI21x1_ASAP7_75t_R _11076_ (.A1(_04946_),
    .A2(_04964_),
    .B(_04987_),
    .Y(_04988_));
 NAND2x1_ASAP7_75t_R _11077_ (.A(net3304),
    .B(_04988_),
    .Y(_04989_));
 XOR2x2_ASAP7_75t_R _11078_ (.A(_04973_),
    .B(net3327),
    .Y(_04990_));
 AOI21x1_ASAP7_75t_R _11079_ (.A1(_04982_),
    .A2(_04989_),
    .B(_04990_),
    .Y(_04991_));
 NAND2x1_ASAP7_75t_R _11080_ (.A(net3261),
    .B(_04991_),
    .Y(_04992_));
 XOR2x2_ASAP7_75t_R _11081_ (.A(_04965_),
    .B(net4198),
    .Y(_04993_));
 INVx1_ASAP7_75t_R _11082_ (.A(_04978_),
    .Y(_04994_));
 OAI21x1_ASAP7_75t_R _11083_ (.A1(_04953_),
    .A2(_04963_),
    .B(net3305),
    .Y(_04995_));
 OAI21x1_ASAP7_75t_R _11084_ (.A1(_04976_),
    .A2(_04994_),
    .B(_04995_),
    .Y(_04996_));
 NOR2x1_ASAP7_75t_R _11085_ (.A(_04953_),
    .B(_04963_),
    .Y(_04997_));
 NAND2x1_ASAP7_75t_R _11086_ (.A(net3370),
    .B(net3306),
    .Y(_04998_));
 AOI21x1_ASAP7_75t_R _11087_ (.A1(net3311),
    .A2(_04998_),
    .B(net3309),
    .Y(_04999_));
 AOI21x1_ASAP7_75t_R _11088_ (.A1(net3287),
    .A2(_04997_),
    .B(_04999_),
    .Y(_05000_));
 NAND2x1_ASAP7_75t_R _11089_ (.A(_04996_),
    .B(_05000_),
    .Y(_05001_));
 INVx1_ASAP7_75t_R _11090_ (.A(_04983_),
    .Y(_05002_));
 AOI211x1_ASAP7_75t_R _11091_ (.A1(_04964_),
    .A2(_04946_),
    .B(_05002_),
    .C(_04987_),
    .Y(_05003_));
 XOR2x2_ASAP7_75t_R _11092_ (.A(_04973_),
    .B(net3326),
    .Y(_05004_));
 OAI21x1_ASAP7_75t_R _11093_ (.A1(_05001_),
    .A2(_05003_),
    .B(_05004_),
    .Y(_05005_));
 NAND2x1_ASAP7_75t_R _11094_ (.A(_04993_),
    .B(_05005_),
    .Y(_05006_));
 NAND2x2_ASAP7_75t_R _11095_ (.A(_04992_),
    .B(_05006_),
    .Y(_05007_));
 INVx2_ASAP7_75t_R _11096_ (.A(_05007_),
    .Y(_05008_));
 OR3x1_ASAP7_75t_R _11097_ (.A(net4415),
    .B(net4416),
    .C(net4357),
    .Y(_05009_));
 XOR2x2_ASAP7_75t_R _11098_ (.A(_05009_),
    .B(net4413),
    .Y(_05010_));
 INVx1_ASAP7_75t_R _11099_ (.A(_05010_),
    .Y(_05011_));
 NOR2x1_ASAP7_75t_R _11100_ (.A(net4118),
    .B(_05005_),
    .Y(_05012_));
 NOR2x1_ASAP7_75t_R _11101_ (.A(net4198),
    .B(_04991_),
    .Y(_05013_));
 OA21x2_ASAP7_75t_R _11102_ (.A1(_05012_),
    .A2(_05013_),
    .B(net3261),
    .Y(_05014_));
 OAI21x1_ASAP7_75t_R _11103_ (.A1(_04990_),
    .A2(_04982_),
    .B(_04989_),
    .Y(_05015_));
 XOR2x2_ASAP7_75t_R _11104_ (.A(_05015_),
    .B(net3256),
    .Y(_05016_));
 XOR2x2_ASAP7_75t_R _11105_ (.A(_04983_),
    .B(net4119),
    .Y(_05017_));
 OAI21x1_ASAP7_75t_R _11106_ (.A1(_04953_),
    .A2(_04963_),
    .B(net3304),
    .Y(_05018_));
 OAI21x1_ASAP7_75t_R _11107_ (.A1(net3271),
    .A2(_05017_),
    .B(_05018_),
    .Y(_05019_));
 NAND2x1_ASAP7_75t_R _11108_ (.A(net3252),
    .B(_04991_),
    .Y(_05020_));
 XOR2x2_ASAP7_75t_R _11109_ (.A(net3257),
    .B(_05019_),
    .Y(_05021_));
 NAND2x1_ASAP7_75t_R _11110_ (.A(_05021_),
    .B(_05005_),
    .Y(_05022_));
 NAND2x1_ASAP7_75t_R _11111_ (.A(_05020_),
    .B(_05022_),
    .Y(_05023_));
 NOR2x1_ASAP7_75t_R _11112_ (.A(_05016_),
    .B(_05023_),
    .Y(_05024_));
 NAND2x1_ASAP7_75t_R _11113_ (.A(_05014_),
    .B(_05024_),
    .Y(_05025_));
 NAND2x1_ASAP7_75t_R _11114_ (.A(net4118),
    .B(_05005_),
    .Y(_05026_));
 NAND2x1_ASAP7_75t_R _11115_ (.A(net4198),
    .B(_04991_),
    .Y(_05027_));
 INVx1_ASAP7_75t_R _11116_ (.A(net3261),
    .Y(_05028_));
 AO21x1_ASAP7_75t_R _11117_ (.A1(_05026_),
    .A2(_05027_),
    .B(_05028_),
    .Y(_05029_));
 AOI21x1_ASAP7_75t_R _11118_ (.A1(net3253),
    .A2(net3241),
    .B(net3254),
    .Y(_05030_));
 NAND2x1_ASAP7_75t_R _11119_ (.A(net3256),
    .B(_05030_),
    .Y(_05031_));
 XOR2x2_ASAP7_75t_R _11120_ (.A(_05031_),
    .B(net3260),
    .Y(_05032_));
 AOI21x1_ASAP7_75t_R _11121_ (.A1(_05029_),
    .A2(_05024_),
    .B(_05032_),
    .Y(_05033_));
 OAI21x1_ASAP7_75t_R _11122_ (.A1(net4197),
    .A2(_05025_),
    .B(_05033_),
    .Y(_05034_));
 AND3x1_ASAP7_75t_R _11123_ (.A(_04990_),
    .B(net3304),
    .C(net3258),
    .Y(_05035_));
 AOI21x1_ASAP7_75t_R _11124_ (.A1(net3258),
    .A2(net3230),
    .B(net3252),
    .Y(_05036_));
 XOR2x2_ASAP7_75t_R _11125_ (.A(_05015_),
    .B(net3259),
    .Y(_05037_));
 OAI21x1_ASAP7_75t_R _11126_ (.A1(_05035_),
    .A2(_05036_),
    .B(_05037_),
    .Y(_05038_));
 XOR2x2_ASAP7_75t_R _11127_ (.A(_05031_),
    .B(net3255),
    .Y(_05039_));
 OAI21x1_ASAP7_75t_R _11128_ (.A1(_05007_),
    .A2(_05038_),
    .B(_05039_),
    .Y(_05040_));
 INVx1_ASAP7_75t_R _11129_ (.A(_05023_),
    .Y(_05041_));
 NAND2x1_ASAP7_75t_R _11130_ (.A(_05007_),
    .B(_05041_),
    .Y(_05042_));
 NAND2x1_ASAP7_75t_R _11131_ (.A(net3256),
    .B(net3229),
    .Y(_05043_));
 NAND2x1_ASAP7_75t_R _11132_ (.A(net3259),
    .B(net3228),
    .Y(_05044_));
 AOI21x1_ASAP7_75t_R _11133_ (.A1(_05043_),
    .A2(_05044_),
    .B(net3255),
    .Y(_05045_));
 OAI21x1_ASAP7_75t_R _11134_ (.A1(_05013_),
    .A2(_05012_),
    .B(_05011_),
    .Y(_05046_));
 NAND2x1_ASAP7_75t_R _11135_ (.A(_05045_),
    .B(_05046_),
    .Y(_05047_));
 NOR2x1_ASAP7_75t_R _11136_ (.A(_05042_),
    .B(_05047_),
    .Y(_05048_));
 XOR2x2_ASAP7_75t_R _11137_ (.A(_05046_),
    .B(_05008_),
    .Y(_05049_));
 OAI21x1_ASAP7_75t_R _11138_ (.A1(_05040_),
    .A2(_05048_),
    .B(_05049_),
    .Y(_05050_));
 OAI21x1_ASAP7_75t_R _11139_ (.A1(net3188),
    .A2(_05034_),
    .B(_05050_),
    .Y(_05051_));
 OA21x2_ASAP7_75t_R _11140_ (.A1(_05046_),
    .A2(net3240),
    .B(_05041_),
    .Y(_05052_));
 AOI21x1_ASAP7_75t_R _11141_ (.A1(_05032_),
    .A2(_05052_),
    .B(net3214),
    .Y(_05053_));
 AO21x1_ASAP7_75t_R _11142_ (.A1(net3214),
    .A2(_05052_),
    .B(_05053_),
    .Y(_05054_));
 INVx1_ASAP7_75t_R _11143_ (.A(_05054_),
    .Y(_05055_));
 OAI22x1_ASAP7_75t_R _11144_ (.A1(_05024_),
    .A2(_05032_),
    .B1(net4262),
    .B2(_05029_),
    .Y(_05056_));
 XOR2x2_ASAP7_75t_R _11145_ (.A(_05056_),
    .B(net3187),
    .Y(_05057_));
 NOR2x1_ASAP7_75t_R _11146_ (.A(_05057_),
    .B(_05051_),
    .Y(_05058_));
 NOR2x1_ASAP7_75t_R _11147_ (.A(net4414),
    .B(net4320),
    .Y(_05059_));
 XOR2x2_ASAP7_75t_R _11148_ (.A(_05059_),
    .B(net4514),
    .Y(_05060_));
 NAND2x1_ASAP7_75t_R _11149_ (.A(net4197),
    .B(_05033_),
    .Y(_05061_));
 NOR2x1_ASAP7_75t_R _11150_ (.A(_05029_),
    .B(_05038_),
    .Y(_05062_));
 OAI21x1_ASAP7_75t_R _11151_ (.A1(_05014_),
    .A2(_05038_),
    .B(_05039_),
    .Y(_05063_));
 OAI21x1_ASAP7_75t_R _11152_ (.A1(_05062_),
    .A2(_05063_),
    .B(net4262),
    .Y(_05064_));
 NAND2x1_ASAP7_75t_R _11153_ (.A(net3215),
    .B(net3216),
    .Y(_05065_));
 INVx1_ASAP7_75t_R _11154_ (.A(_05065_),
    .Y(_05066_));
 AOI21x1_ASAP7_75t_R _11155_ (.A1(_05061_),
    .A2(_05064_),
    .B(_05066_),
    .Y(_05067_));
 NAND2x1_ASAP7_75t_R _11156_ (.A(_05060_),
    .B(_05067_),
    .Y(_05068_));
 OAI21x1_ASAP7_75t_R _11157_ (.A1(net3138),
    .A2(net3124),
    .B(net3137),
    .Y(_05069_));
 NOR2x1_ASAP7_75t_R _11158_ (.A(net3139),
    .B(_05069_),
    .Y(_05070_));
 XOR2x2_ASAP7_75t_R _11159_ (.A(_05056_),
    .B(net3200),
    .Y(_05071_));
 INVx1_ASAP7_75t_R _11160_ (.A(_05060_),
    .Y(_05072_));
 NOR2x1_ASAP7_75t_R _11161_ (.A(net4262),
    .B(_05063_),
    .Y(_05073_));
 AOI21x1_ASAP7_75t_R _11162_ (.A1(_05025_),
    .A2(_05033_),
    .B(net4197),
    .Y(_05074_));
 OAI21x1_ASAP7_75t_R _11163_ (.A1(_05073_),
    .A2(_05074_),
    .B(net3198),
    .Y(_05075_));
 NOR2x1_ASAP7_75t_R _11164_ (.A(_05072_),
    .B(_05075_),
    .Y(_05076_));
 INVx1_ASAP7_75t_R _11165_ (.A(_05040_),
    .Y(_05077_));
 OAI21x1_ASAP7_75t_R _11166_ (.A1(net3199),
    .A2(_05077_),
    .B(net3188),
    .Y(_05078_));
 INVx1_ASAP7_75t_R _11167_ (.A(net3199),
    .Y(_05079_));
 NAND3x1_ASAP7_75t_R _11168_ (.A(_05040_),
    .B(net3201),
    .C(_05079_),
    .Y(_05080_));
 NAND2x1_ASAP7_75t_R _11169_ (.A(_05078_),
    .B(_05080_),
    .Y(_05081_));
 NAND2x1_ASAP7_75t_R _11170_ (.A(_05071_),
    .B(_05081_),
    .Y(_05082_));
 NOR2x1_ASAP7_75t_R _11171_ (.A(net3136),
    .B(net3135),
    .Y(_05083_));
 INVx1_ASAP7_75t_R _11172_ (.A(_05083_),
    .Y(_05084_));
 OA21x2_ASAP7_75t_R _11173_ (.A1(_05070_),
    .A2(_05071_),
    .B(_05084_),
    .Y(_05085_));
 BUFx3_ASAP7_75t_R place2952 (.A(_02269_),
    .Y(net2952));
 XOR2x2_ASAP7_75t_R _11175_ (.A(_05069_),
    .B(net3151),
    .Y(_05087_));
 AOI21x1_ASAP7_75t_R _11176_ (.A1(_05068_),
    .A2(_05058_),
    .B(_05055_),
    .Y(_05088_));
 OAI21x1_ASAP7_75t_R _11177_ (.A1(_05073_),
    .A2(_05074_),
    .B(net4196),
    .Y(_05089_));
 NAND2x1_ASAP7_75t_R _11178_ (.A(net3186),
    .B(_05040_),
    .Y(_05090_));
 AO21x1_ASAP7_75t_R _11179_ (.A1(_05063_),
    .A2(net4197),
    .B(_05065_),
    .Y(_05091_));
 NAND2x1_ASAP7_75t_R _11180_ (.A(_05090_),
    .B(_05091_),
    .Y(_05092_));
 XNOR2x2_ASAP7_75t_R _11181_ (.A(_05089_),
    .B(_05092_),
    .Y(_05093_));
 INVx1_ASAP7_75t_R _11182_ (.A(net3163),
    .Y(_05094_));
 NAND2x1_ASAP7_75t_R _11183_ (.A(_05094_),
    .B(_05088_),
    .Y(_05095_));
 OAI21x1_ASAP7_75t_R _11184_ (.A1(_05088_),
    .A2(_05093_),
    .B(_05095_),
    .Y(_05096_));
 NOR2x2_ASAP7_75t_R _11185_ (.A(_05087_),
    .B(_05096_),
    .Y(_05097_));
 BUFx3_ASAP7_75t_R place2951 (.A(_02283_),
    .Y(net2951));
 NOR2x1_ASAP7_75t_R _11187_ (.A(net4407),
    .B(net4320),
    .Y(_05099_));
 XOR2x2_ASAP7_75t_R _11188_ (.A(_05099_),
    .B(net4517),
    .Y(_05100_));
 NAND2x1_ASAP7_75t_R _11189_ (.A(net4195),
    .B(_05088_),
    .Y(_05101_));
 OAI21x1_ASAP7_75t_R _11190_ (.A1(_05076_),
    .A2(_05082_),
    .B(net3152),
    .Y(_05102_));
 NAND2x1_ASAP7_75t_R _11191_ (.A(net4117),
    .B(_05102_),
    .Y(_05103_));
 NAND2x1_ASAP7_75t_R _11192_ (.A(net3164),
    .B(net3178),
    .Y(_05104_));
 INVx1_ASAP7_75t_R _11193_ (.A(net3149),
    .Y(_05105_));
 AOI21x1_ASAP7_75t_R _11194_ (.A1(_05101_),
    .A2(_05103_),
    .B(_05105_),
    .Y(_05106_));
 NAND2x1_ASAP7_75t_R _11195_ (.A(net4194),
    .B(_05106_),
    .Y(_05107_));
 OAI21x1_ASAP7_75t_R _11196_ (.A1(net3095),
    .A2(_05097_),
    .B(_05107_),
    .Y(_05108_));
 NOR2x1_ASAP7_75t_R _11197_ (.A(_05093_),
    .B(_05088_),
    .Y(_05109_));
 NOR2x1_ASAP7_75t_R _11198_ (.A(net3163),
    .B(_05102_),
    .Y(_05110_));
 NOR2x1_ASAP7_75t_R _11199_ (.A(_05109_),
    .B(_05110_),
    .Y(_05111_));
 XOR2x2_ASAP7_75t_R _11200_ (.A(_05108_),
    .B(net3092),
    .Y(_05112_));
 NAND2x1_ASAP7_75t_R _11201_ (.A(net3150),
    .B(_05088_),
    .Y(_05113_));
 XOR2x2_ASAP7_75t_R _11202_ (.A(_05104_),
    .B(net4117),
    .Y(_05114_));
 AO21x1_ASAP7_75t_R _11203_ (.A1(_05084_),
    .A2(net3152),
    .B(_05114_),
    .Y(_05115_));
 NAND2x1_ASAP7_75t_R _11204_ (.A(_05113_),
    .B(_05115_),
    .Y(_05116_));
 INVx1_ASAP7_75t_R _11205_ (.A(_05116_),
    .Y(_05117_));
 XOR2x2_ASAP7_75t_R _11206_ (.A(_05069_),
    .B(net3139),
    .Y(_05118_));
 NAND2x1_ASAP7_75t_R _11207_ (.A(_05118_),
    .B(_05111_),
    .Y(_05119_));
 NOR2x1_ASAP7_75t_R _11208_ (.A(_05116_),
    .B(_05119_),
    .Y(_05120_));
 INVx1_ASAP7_75t_R _11209_ (.A(_05100_),
    .Y(_05121_));
 NOR2x2_ASAP7_75t_R _11210_ (.A(net4195),
    .B(_05088_),
    .Y(_05122_));
 NOR2x1_ASAP7_75t_R _11211_ (.A(net4117),
    .B(_05102_),
    .Y(_05123_));
 NOR2x1_ASAP7_75t_R _11212_ (.A(net3100),
    .B(_05123_),
    .Y(_05124_));
 NOR2x1_ASAP7_75t_R _11213_ (.A(_05121_),
    .B(_05124_),
    .Y(_05125_));
 OAI21x1_ASAP7_75t_R _11214_ (.A1(_05085_),
    .A2(_05120_),
    .B(net3077),
    .Y(_05126_));
 AND3x1_ASAP7_75t_R _11215_ (.A(_05125_),
    .B(_05085_),
    .C(net3149),
    .Y(_05127_));
 AOI21x1_ASAP7_75t_R _11216_ (.A1(_05117_),
    .A2(_05126_),
    .B(_05127_),
    .Y(_05128_));
 NOR2x1_ASAP7_75t_R _11217_ (.A(_05112_),
    .B(_05128_),
    .Y(_05129_));
 OAI21x1_ASAP7_75t_R _11218_ (.A1(_05122_),
    .A2(_05123_),
    .B(net3149),
    .Y(_05130_));
 NOR2x1_ASAP7_75t_R _11219_ (.A(_05121_),
    .B(_05130_),
    .Y(_05131_));
 NOR2x1_ASAP7_75t_R _11220_ (.A(net3093),
    .B(_05131_),
    .Y(_05132_));
 INVx1_ASAP7_75t_R _11221_ (.A(_05085_),
    .Y(_05133_));
 OAI21x1_ASAP7_75t_R _11222_ (.A1(_05119_),
    .A2(_05131_),
    .B(_05133_),
    .Y(_05134_));
 NAND2x1_ASAP7_75t_R _11223_ (.A(_05132_),
    .B(_05134_),
    .Y(_05135_));
 XOR2x2_ASAP7_75t_R _11224_ (.A(_05135_),
    .B(net3102),
    .Y(_05136_));
 AO21x1_ASAP7_75t_R _11225_ (.A1(net4515),
    .A2(net4457),
    .B(net4320),
    .Y(_05137_));
 XNOR2x2_ASAP7_75t_R _11226_ (.A(net4611),
    .B(_05137_),
    .Y(_05138_));
 INVx1_ASAP7_75t_R _11227_ (.A(_05138_),
    .Y(_05139_));
 OA21x2_ASAP7_75t_R _11228_ (.A1(net3022),
    .A2(net3036),
    .B(net4115),
    .Y(_05140_));
 INVx1_ASAP7_75t_R _11229_ (.A(_05140_),
    .Y(_05141_));
 INVx1_ASAP7_75t_R _11230_ (.A(net3091),
    .Y(_05142_));
 AOI21x1_ASAP7_75t_R _11231_ (.A1(_05097_),
    .A2(_05107_),
    .B(_05085_),
    .Y(_05143_));
 NAND2x1_ASAP7_75t_R _11232_ (.A(net4194),
    .B(_05143_),
    .Y(_05144_));
 NAND2x1_ASAP7_75t_R _11233_ (.A(net4116),
    .B(_05134_),
    .Y(_05145_));
 AOI21x1_ASAP7_75t_R _11234_ (.A1(_05144_),
    .A2(_05145_),
    .B(_05139_),
    .Y(_05146_));
 NAND2x1_ASAP7_75t_R _11235_ (.A(net3076),
    .B(_05146_),
    .Y(_05147_));
 AOI21x1_ASAP7_75t_R _11236_ (.A1(_05129_),
    .A2(_05147_),
    .B(_05136_),
    .Y(_05148_));
 NAND2x1_ASAP7_75t_R _11237_ (.A(net4193),
    .B(_05148_),
    .Y(_05149_));
 NAND2x1_ASAP7_75t_R _11238_ (.A(_05141_),
    .B(_05149_),
    .Y(_05150_));
 INVx1_ASAP7_75t_R _11239_ (.A(_05150_),
    .Y(_05151_));
 AO21x1_ASAP7_75t_R _11240_ (.A1(_05146_),
    .A2(net3076),
    .B(net3037),
    .Y(_05152_));
 XOR2x2_ASAP7_75t_R _11241_ (.A(_05135_),
    .B(net3101),
    .Y(_05153_));
 AOI211x1_ASAP7_75t_R _11242_ (.A1(net3078),
    .A2(net3090),
    .B(net3094),
    .C(net4116),
    .Y(_05154_));
 NOR2x1_ASAP7_75t_R _11243_ (.A(net4194),
    .B(net3062),
    .Y(_05155_));
 OAI21x1_ASAP7_75t_R _11244_ (.A1(_05154_),
    .A2(_05155_),
    .B(net3076),
    .Y(_05156_));
 NOR2x1_ASAP7_75t_R _11245_ (.A(net4115),
    .B(_05156_),
    .Y(_05157_));
 OAI21x1_ASAP7_75t_R _11246_ (.A1(_05153_),
    .A2(_05157_),
    .B(net3037),
    .Y(_05158_));
 OAI21x1_ASAP7_75t_R _11247_ (.A1(_05152_),
    .A2(_05148_),
    .B(_05158_),
    .Y(_05159_));
 INVx2_ASAP7_75t_R _11248_ (.A(_05159_),
    .Y(_05160_));
 OAI21x1_ASAP7_75t_R _11249_ (.A1(_05154_),
    .A2(_05155_),
    .B(net4193),
    .Y(_05161_));
 XOR2x2_ASAP7_75t_R _11250_ (.A(net3091),
    .B(net4194),
    .Y(_05162_));
 NAND2x1_ASAP7_75t_R _11251_ (.A(_05142_),
    .B(net3062),
    .Y(_05163_));
 OAI21x1_ASAP7_75t_R _11252_ (.A1(net3062),
    .A2(_05162_),
    .B(_05163_),
    .Y(_05164_));
 INVx1_ASAP7_75t_R _11253_ (.A(net3033),
    .Y(_05165_));
 AOI211x1_ASAP7_75t_R _11254_ (.A1(net3022),
    .A2(net3034),
    .B(_05165_),
    .C(net3036),
    .Y(_05166_));
 XOR2x2_ASAP7_75t_R _11255_ (.A(_05161_),
    .B(_05164_),
    .Y(_05167_));
 NOR2x2_ASAP7_75t_R _11256_ (.A(_05167_),
    .B(_05148_),
    .Y(_05168_));
 NOR2x2_ASAP7_75t_R _11257_ (.A(_05166_),
    .B(_05168_),
    .Y(_05169_));
 NAND2x2_ASAP7_75t_R _11258_ (.A(_05160_),
    .B(_05169_),
    .Y(_05170_));
 OR3x1_ASAP7_75t_R _11259_ (.A(net4415),
    .B(net4416),
    .C(_04440_),
    .Y(_05171_));
 XNOR2x2_ASAP7_75t_R _11260_ (.A(net4516),
    .B(_05171_),
    .Y(_05172_));
 INVx1_ASAP7_75t_R _11261_ (.A(_05172_),
    .Y(_05173_));
 AOI211x1_ASAP7_75t_R _11262_ (.A1(net3022),
    .A2(_05156_),
    .B(net3036),
    .C(net4115),
    .Y(_05174_));
 NAND2x1_ASAP7_75t_R _11263_ (.A(net3046),
    .B(net3045),
    .Y(_05175_));
 OAI21x1_ASAP7_75t_R _11264_ (.A1(_05140_),
    .A2(_05174_),
    .B(_05175_),
    .Y(_05176_));
 NOR2x1_ASAP7_75t_R _11265_ (.A(_05173_),
    .B(_05176_),
    .Y(_05177_));
 INVx1_ASAP7_75t_R _11266_ (.A(net3047),
    .Y(_05178_));
 NAND2x1_ASAP7_75t_R _11267_ (.A(_05178_),
    .B(_05153_),
    .Y(_05179_));
 AOI21x1_ASAP7_75t_R _11268_ (.A1(_05153_),
    .A2(_05179_),
    .B(_05152_),
    .Y(_05180_));
 XOR2x2_ASAP7_75t_R _11269_ (.A(_05180_),
    .B(net3032),
    .Y(_05181_));
 INVx2_ASAP7_75t_R _11270_ (.A(_05181_),
    .Y(_05182_));
 OAI21x1_ASAP7_75t_R _11271_ (.A1(_05170_),
    .A2(_05177_),
    .B(_05182_),
    .Y(_05183_));
 NOR2x1_ASAP7_75t_R _11272_ (.A(net4313),
    .B(net2976),
    .Y(_05184_));
 NOR2x1_ASAP7_75t_R _11273_ (.A(net4260),
    .B(net2993),
    .Y(_05185_));
 OAI21x1_ASAP7_75t_R _11274_ (.A1(_05184_),
    .A2(_05185_),
    .B(net2962),
    .Y(_05186_));
 OAI21x1_ASAP7_75t_R _11275_ (.A1(net2977),
    .A2(net2963),
    .B(_05186_),
    .Y(_05187_));
 NOR2x1_ASAP7_75t_R _11276_ (.A(net4260),
    .B(_05151_),
    .Y(_05188_));
 NOR2x1_ASAP7_75t_R _11277_ (.A(net4115),
    .B(net3013),
    .Y(_05189_));
 INVx1_ASAP7_75t_R _11278_ (.A(_05175_),
    .Y(_05190_));
 XOR2x2_ASAP7_75t_R _11279_ (.A(_05189_),
    .B(_05190_),
    .Y(_05191_));
 INVx1_ASAP7_75t_R _11280_ (.A(_05191_),
    .Y(_05192_));
 AOI21x1_ASAP7_75t_R _11281_ (.A1(_05188_),
    .A2(_05183_),
    .B(_05192_),
    .Y(_05193_));
 NAND2x1_ASAP7_75t_R _11282_ (.A(net2990),
    .B(_05183_),
    .Y(_05194_));
 INVx1_ASAP7_75t_R _11283_ (.A(_05194_),
    .Y(_05195_));
 INVx1_ASAP7_75t_R _11284_ (.A(net2990),
    .Y(_05196_));
 AOI21x1_ASAP7_75t_R _11285_ (.A1(net2998),
    .A2(_05196_),
    .B(net2991),
    .Y(_05197_));
 OAI21x1_ASAP7_75t_R _11286_ (.A1(net4259),
    .A2(net2999),
    .B(_05169_),
    .Y(_05198_));
 AOI21x1_ASAP7_75t_R _11287_ (.A1(_05182_),
    .A2(net3000),
    .B(_05198_),
    .Y(_05199_));
 NOR2x1_ASAP7_75t_R _11288_ (.A(_05197_),
    .B(_05199_),
    .Y(_05200_));
 OAI21x1_ASAP7_75t_R _11289_ (.A1(_05193_),
    .A2(_05195_),
    .B(_05200_),
    .Y(_05201_));
 XOR2x2_ASAP7_75t_R _11290_ (.A(_05199_),
    .B(net2992),
    .Y(_05202_));
 INVx2_ASAP7_75t_R _11291_ (.A(_05202_),
    .Y(_05203_));
 OAI21x1_ASAP7_75t_R _11292_ (.A1(_05187_),
    .A2(_05201_),
    .B(_05203_),
    .Y(_05204_));
 NAND3x1_ASAP7_75t_R _11293_ (.A(net2999),
    .B(net2991),
    .C(net2992),
    .Y(_05205_));
 NAND3x1_ASAP7_75t_R _11294_ (.A(_05205_),
    .B(net4313),
    .C(net2989),
    .Y(_05206_));
 AO21x1_ASAP7_75t_R _11295_ (.A1(_05182_),
    .A2(_05170_),
    .B(net4313),
    .Y(_05207_));
 NOR2x1_ASAP7_75t_R _11296_ (.A(net4515),
    .B(net4320),
    .Y(_05208_));
 XOR2x2_ASAP7_75t_R _11297_ (.A(_05208_),
    .B(net4553),
    .Y(_05209_));
 INVx1_ASAP7_75t_R _11298_ (.A(_05209_),
    .Y(_05210_));
 AO21x1_ASAP7_75t_R _11299_ (.A1(_05206_),
    .A2(_05207_),
    .B(_05210_),
    .Y(_05211_));
 INVx1_ASAP7_75t_R _11300_ (.A(_05211_),
    .Y(_05212_));
 AO21x1_ASAP7_75t_R _11301_ (.A1(_05204_),
    .A2(_05212_),
    .B(net2932),
    .Y(_05213_));
 NAND3x1_ASAP7_75t_R _11302_ (.A(_05204_),
    .B(_05212_),
    .C(net2932),
    .Y(_05214_));
 INVx1_ASAP7_75t_R _11303_ (.A(_05207_),
    .Y(_05215_));
 NOR2x1_ASAP7_75t_R _11304_ (.A(net4261),
    .B(net2962),
    .Y(_05216_));
 OAI21x1_ASAP7_75t_R _11305_ (.A1(_05215_),
    .A2(_05216_),
    .B(net2993),
    .Y(_05217_));
 NOR2x1_ASAP7_75t_R _11306_ (.A(net4113),
    .B(_05217_),
    .Y(_05218_));
 NOR2x1_ASAP7_75t_R _11307_ (.A(_05193_),
    .B(_05195_),
    .Y(_05219_));
 OAI21x1_ASAP7_75t_R _11308_ (.A1(_05203_),
    .A2(_05218_),
    .B(net2919),
    .Y(_05220_));
 AOI21x1_ASAP7_75t_R _11309_ (.A1(_05207_),
    .A2(_05206_),
    .B(net2977),
    .Y(_05221_));
 AOI21x1_ASAP7_75t_R _11310_ (.A1(net4192),
    .A2(_05221_),
    .B(_05219_),
    .Y(_05222_));
 OAI21x1_ASAP7_75t_R _11311_ (.A1(net2944),
    .A2(net2942),
    .B(_05222_),
    .Y(_05223_));
 NAND2x1_ASAP7_75t_R _11312_ (.A(_05220_),
    .B(_05223_),
    .Y(_05224_));
 AOI21x1_ASAP7_75t_R _11313_ (.A1(_05213_),
    .A2(_05214_),
    .B(_05224_),
    .Y(_05225_));
 INVx1_ASAP7_75t_R _11314_ (.A(_05188_),
    .Y(_05226_));
 NAND2x1_ASAP7_75t_R _11315_ (.A(net3033),
    .B(net3012),
    .Y(_05227_));
 INVx1_ASAP7_75t_R _11316_ (.A(_05167_),
    .Y(_05228_));
 INVx1_ASAP7_75t_R _11317_ (.A(net3022),
    .Y(_05229_));
 OAI21x1_ASAP7_75t_R _11318_ (.A1(net3021),
    .A2(_05229_),
    .B(net3035),
    .Y(_05230_));
 NAND2x1_ASAP7_75t_R _11319_ (.A(_05228_),
    .B(_05230_),
    .Y(_05231_));
 NAND2x1_ASAP7_75t_R _11320_ (.A(_05227_),
    .B(_05231_),
    .Y(_05232_));
 NOR2x1_ASAP7_75t_R _11321_ (.A(net3000),
    .B(_05232_),
    .Y(_05233_));
 AOI21x1_ASAP7_75t_R _11322_ (.A1(net2987),
    .A2(_05233_),
    .B(net2998),
    .Y(_05234_));
 OAI21x1_ASAP7_75t_R _11323_ (.A1(_05226_),
    .A2(_05234_),
    .B(net2987),
    .Y(_05235_));
 OAI21x1_ASAP7_75t_R _11324_ (.A1(net2990),
    .A2(net2988),
    .B(_05232_),
    .Y(_05236_));
 AOI21x1_ASAP7_75t_R _11325_ (.A1(_05141_),
    .A2(_05149_),
    .B(net3020),
    .Y(_05237_));
 AOI21x1_ASAP7_75t_R _11326_ (.A1(net4313),
    .A2(_05237_),
    .B(_05232_),
    .Y(_05238_));
 OAI21x1_ASAP7_75t_R _11327_ (.A1(net2998),
    .A2(net2992),
    .B(_05238_),
    .Y(_05239_));
 NAND2x1_ASAP7_75t_R _11328_ (.A(_05236_),
    .B(_05239_),
    .Y(_05240_));
 AOI21x1_ASAP7_75t_R _11329_ (.A1(_05235_),
    .A2(net2945),
    .B(_05240_),
    .Y(_05241_));
 AOI211x1_ASAP7_75t_R _11330_ (.A1(_05241_),
    .A2(_05217_),
    .B(net2942),
    .C(net4113),
    .Y(_05242_));
 OAI21x1_ASAP7_75t_R _11331_ (.A1(net4113),
    .A2(_05217_),
    .B(_05241_),
    .Y(_05243_));
 AOI21x1_ASAP7_75t_R _11332_ (.A1(net2930),
    .A2(_05243_),
    .B(net4192),
    .Y(_05244_));
 NAND2x1_ASAP7_75t_R _11333_ (.A(net2960),
    .B(net2961),
    .Y(_05245_));
 OAI21x1_ASAP7_75t_R _11334_ (.A1(_05242_),
    .A2(_05244_),
    .B(_05245_),
    .Y(_05246_));
 AOI21x1_ASAP7_75t_R _11335_ (.A1(net4192),
    .A2(_05221_),
    .B(_05201_),
    .Y(_05247_));
 AO21x1_ASAP7_75t_R _11336_ (.A1(_05223_),
    .A2(net2929),
    .B(_05247_),
    .Y(_05248_));
 BUFx3_ASAP7_75t_R place2957 (.A(_06317_),
    .Y(net2957));
 INVx3_ASAP7_75t_R _11338_ (.A(_05248_),
    .Y(_05250_));
 OR3x1_ASAP7_75t_R _11339_ (.A(net4415),
    .B(net4416),
    .C(_04438_),
    .Y(_05251_));
 XOR2x2_ASAP7_75t_R _11340_ (.A(_05251_),
    .B(net4610),
    .Y(_05252_));
 INVx1_ASAP7_75t_R _11341_ (.A(_05252_),
    .Y(_05253_));
 AOI211x1_ASAP7_75t_R _11342_ (.A1(_05225_),
    .A2(_05246_),
    .B(_05250_),
    .C(_05253_),
    .Y(_05254_));
 OAI21x1_ASAP7_75t_R _11343_ (.A1(net4257),
    .A2(net2871),
    .B(_05225_),
    .Y(_05255_));
 AOI21x1_ASAP7_75t_R _11344_ (.A1(net2870),
    .A2(_05255_),
    .B(net4312),
    .Y(_05256_));
 NOR2x1_ASAP7_75t_R _11345_ (.A(net2838),
    .B(_05256_),
    .Y(_05257_));
 NOR2x1_ASAP7_75t_R _11346_ (.A(_04368_),
    .B(_05257_),
    .Y(_05258_));
 NOR2x1_ASAP7_75t_R _11347_ (.A(net4257),
    .B(_05246_),
    .Y(_05259_));
 AOI211x1_ASAP7_75t_R _11348_ (.A1(_05201_),
    .A2(_05203_),
    .B(net2932),
    .C(_05211_),
    .Y(_05260_));
 INVx1_ASAP7_75t_R _11349_ (.A(_05187_),
    .Y(_05261_));
 AOI21x1_ASAP7_75t_R _11350_ (.A1(_05212_),
    .A2(_05204_),
    .B(_05261_),
    .Y(_05262_));
 NOR2x1_ASAP7_75t_R _11351_ (.A(_05260_),
    .B(_05262_),
    .Y(_05263_));
 INVx1_ASAP7_75t_R _11352_ (.A(_05263_),
    .Y(_05264_));
 OAI21x1_ASAP7_75t_R _11353_ (.A1(net2870),
    .A2(_05259_),
    .B(net2852),
    .Y(_05265_));
 INVx1_ASAP7_75t_R _11354_ (.A(_05224_),
    .Y(_05266_));
 OAI21x1_ASAP7_75t_R _11355_ (.A1(net2943),
    .A2(net2900),
    .B(net4114),
    .Y(_05267_));
 INVx1_ASAP7_75t_R _11356_ (.A(_05242_),
    .Y(_05268_));
 AOI21x1_ASAP7_75t_R _11357_ (.A1(_05267_),
    .A2(_05268_),
    .B(_05253_),
    .Y(_05269_));
 AOI21x1_ASAP7_75t_R _11358_ (.A1(net2941),
    .A2(_05269_),
    .B(_05264_),
    .Y(_05270_));
 OAI21x1_ASAP7_75t_R _11359_ (.A1(_05250_),
    .A2(_05266_),
    .B(_05270_),
    .Y(_05271_));
 NAND2x1_ASAP7_75t_R _11360_ (.A(_05265_),
    .B(_05271_),
    .Y(_05272_));
 INVx1_ASAP7_75t_R _11361_ (.A(_05269_),
    .Y(_05273_));
 INVx1_ASAP7_75t_R _11362_ (.A(net2941),
    .Y(_05274_));
 NAND2x1_ASAP7_75t_R _11363_ (.A(net2931),
    .B(net2901),
    .Y(_05275_));
 XOR2x2_ASAP7_75t_R _11364_ (.A(_05245_),
    .B(net4192),
    .Y(_05276_));
 OAI21x1_ASAP7_75t_R _11365_ (.A1(net2943),
    .A2(net2900),
    .B(_05276_),
    .Y(_05277_));
 OAI21x1_ASAP7_75t_R _11366_ (.A1(_05274_),
    .A2(_05275_),
    .B(_05277_),
    .Y(_05278_));
 INVx1_ASAP7_75t_R _11367_ (.A(_05278_),
    .Y(_05279_));
 AOI21x1_ASAP7_75t_R _11368_ (.A1(_05279_),
    .A2(net2855),
    .B(net2854),
    .Y(_05280_));
 NOR2x1_ASAP7_75t_R _11369_ (.A(net2851),
    .B(_05280_),
    .Y(_05281_));
 NAND2x1_ASAP7_75t_R _11370_ (.A(net2869),
    .B(_05266_),
    .Y(_05282_));
 OAI21x1_ASAP7_75t_R _11371_ (.A1(net2837),
    .A2(net2853),
    .B(net2870),
    .Y(_05283_));
 NOR2x1_ASAP7_75t_R _11372_ (.A(net2902),
    .B(net2883),
    .Y(_05284_));
 INVx1_ASAP7_75t_R _11373_ (.A(_05284_),
    .Y(_05285_));
 AOI21x1_ASAP7_75t_R _11374_ (.A1(net4312),
    .A2(_05283_),
    .B(net2850),
    .Y(_05286_));
 OA31x2_ASAP7_75t_R _11375_ (.A1(net4258),
    .A2(net2870),
    .A3(_05284_),
    .B1(_05278_),
    .Y(_05287_));
 AOI211x1_ASAP7_75t_R _11376_ (.A1(_05282_),
    .A2(net2870),
    .B(_05273_),
    .C(net2941),
    .Y(_05288_));
 NOR2x1_ASAP7_75t_R _11377_ (.A(_05287_),
    .B(_05288_),
    .Y(_05289_));
 OAI21x1_ASAP7_75t_R _11378_ (.A1(_05281_),
    .A2(_05286_),
    .B(_05289_),
    .Y(_05290_));
 XOR2x2_ASAP7_75t_R _11379_ (.A(_05271_),
    .B(net2872),
    .Y(_05291_));
 INVx2_ASAP7_75t_R _11380_ (.A(_05291_),
    .Y(_05292_));
 OAI21x1_ASAP7_75t_R _11381_ (.A1(net2813),
    .A2(_05290_),
    .B(_05292_),
    .Y(_05293_));
 NOR2x1_ASAP7_75t_R _11382_ (.A(_05281_),
    .B(_05286_),
    .Y(_05294_));
 AOI21x1_ASAP7_75t_R _11383_ (.A1(_05258_),
    .A2(_05293_),
    .B(_05294_),
    .Y(_05295_));
 AND3x1_ASAP7_75t_R _11384_ (.A(_05258_),
    .B(net2850),
    .C(_05291_),
    .Y(_05296_));
 OAI21x1_ASAP7_75t_R _11385_ (.A1(_05254_),
    .A2(_05256_),
    .B(_05285_),
    .Y(_05297_));
 INVx1_ASAP7_75t_R _11386_ (.A(_05297_),
    .Y(_05298_));
 NAND2x1_ASAP7_75t_R _11387_ (.A(net4268),
    .B(_05298_),
    .Y(_05299_));
 AOI21x1_ASAP7_75t_R _11388_ (.A1(_05291_),
    .A2(_05299_),
    .B(net2812),
    .Y(_05300_));
 OAI21x1_ASAP7_75t_R _11389_ (.A1(_04368_),
    .A2(_05297_),
    .B(_05289_),
    .Y(_05301_));
 AOI21x1_ASAP7_75t_R _11390_ (.A1(_05292_),
    .A2(net2813),
    .B(_05301_),
    .Y(_05302_));
 NOR2x2_ASAP7_75t_R _11391_ (.A(_05300_),
    .B(_05302_),
    .Y(_05303_));
 OAI21x1_ASAP7_75t_R _11392_ (.A1(_05295_),
    .A2(_05296_),
    .B(_05303_),
    .Y(_05304_));
 OR3x1_ASAP7_75t_R _11393_ (.A(net4415),
    .B(net4416),
    .C(net4608),
    .Y(_05305_));
 XOR2x2_ASAP7_75t_R _11394_ (.A(_05305_),
    .B(net4614),
    .Y(_05306_));
 OR3x1_ASAP7_75t_R _11395_ (.A(_05273_),
    .B(net2928),
    .C(net2870),
    .Y(_05307_));
 OAI21x1_ASAP7_75t_R _11396_ (.A1(net2851),
    .A2(_05280_),
    .B(_05279_),
    .Y(_05308_));
 AOI21x1_ASAP7_75t_R _11397_ (.A1(_05307_),
    .A2(_05308_),
    .B(_05272_),
    .Y(_05309_));
 OA21x2_ASAP7_75t_R _11398_ (.A1(_05309_),
    .A2(_05291_),
    .B(_04368_),
    .Y(_05310_));
 AOI211x1_ASAP7_75t_R _11399_ (.A1(_05309_),
    .A2(_05297_),
    .B(_05291_),
    .C(_04368_),
    .Y(_05311_));
 INVx1_ASAP7_75t_R _11400_ (.A(net2814),
    .Y(_05312_));
 OAI21x1_ASAP7_75t_R _11401_ (.A1(_05310_),
    .A2(_05311_),
    .B(_05312_),
    .Y(_05313_));
 NOR2x1_ASAP7_75t_R _11402_ (.A(_05306_),
    .B(_05313_),
    .Y(_05314_));
 INVx1_ASAP7_75t_R _11403_ (.A(net2813),
    .Y(_05315_));
 INVx1_ASAP7_75t_R _11404_ (.A(_05309_),
    .Y(_05316_));
 NOR2x1_ASAP7_75t_R _11405_ (.A(_04368_),
    .B(net2811),
    .Y(_05317_));
 OAI22x1_ASAP7_75t_R _11406_ (.A1(_05302_),
    .A2(_05315_),
    .B1(_05316_),
    .B2(_05317_),
    .Y(_05318_));
 OAI21x1_ASAP7_75t_R _11407_ (.A1(_05304_),
    .A2(_05314_),
    .B(_05318_),
    .Y(_05319_));
 INVx1_ASAP7_75t_R _11408_ (.A(net2777),
    .Y(_05320_));
 INVx1_ASAP7_75t_R _11409_ (.A(net2785),
    .Y(_05321_));
 AO21x1_ASAP7_75t_R _11410_ (.A1(_05320_),
    .A2(_05321_),
    .B(net2760),
    .Y(_05322_));
 XOR2x2_ASAP7_75t_R _11411_ (.A(_05322_),
    .B(net2761),
    .Y(_05323_));
 NOR2x1_ASAP7_75t_R _11412_ (.A(net2761),
    .B(net2743),
    .Y(_05324_));
 AOI21x1_ASAP7_75t_R _11413_ (.A1(net2743),
    .A2(_05323_),
    .B(_05324_),
    .Y(_05325_));
 INVx1_ASAP7_75t_R _11414_ (.A(_05325_),
    .Y(_05326_));
 AOI21x1_ASAP7_75t_R _11415_ (.A1(_05318_),
    .A2(_05304_),
    .B(net2760),
    .Y(_05327_));
 NOR2x1_ASAP7_75t_R _11416_ (.A(net2785),
    .B(net2777),
    .Y(_05328_));
 XOR2x2_ASAP7_75t_R _11417_ (.A(_05327_),
    .B(_05328_),
    .Y(_05329_));
 OAI21x1_ASAP7_75t_R _11418_ (.A1(_05316_),
    .A2(_05317_),
    .B(net2799),
    .Y(_05330_));
 XOR2x2_ASAP7_75t_R _11419_ (.A(net2814),
    .B(net4207),
    .Y(_05331_));
 NAND2x1_ASAP7_75t_R _11420_ (.A(_05331_),
    .B(_05330_),
    .Y(_05332_));
 OAI21x1_ASAP7_75t_R _11421_ (.A1(net2814),
    .A2(net2773),
    .B(_05332_),
    .Y(_05333_));
 INVx1_ASAP7_75t_R _11422_ (.A(_05333_),
    .Y(_05334_));
 INVx1_ASAP7_75t_R _11423_ (.A(net4311),
    .Y(_05335_));
 OR2x2_ASAP7_75t_R _11424_ (.A(_05310_),
    .B(_05311_),
    .Y(_05336_));
 NAND2x1_ASAP7_75t_R _11425_ (.A(_05335_),
    .B(_05336_),
    .Y(_05337_));
 INVx1_ASAP7_75t_R _11426_ (.A(_05337_),
    .Y(_05338_));
 OAI21x1_ASAP7_75t_R _11427_ (.A1(_05333_),
    .A2(_05304_),
    .B(net2774),
    .Y(_05339_));
 NAND2x1_ASAP7_75t_R _11428_ (.A(_05338_),
    .B(_05339_),
    .Y(_05340_));
 NOR3x1_ASAP7_75t_R _11429_ (.A(net2775),
    .B(net4311),
    .C(net2776),
    .Y(_05341_));
 AOI21x1_ASAP7_75t_R _11430_ (.A1(_05334_),
    .A2(_05340_),
    .B(_05341_),
    .Y(_05342_));
 NAND2x1_ASAP7_75t_R _11431_ (.A(_05329_),
    .B(_05342_),
    .Y(_05343_));
 INVx1_ASAP7_75t_R _11432_ (.A(_05343_),
    .Y(_05344_));
 NOR2x1_ASAP7_75t_R _11433_ (.A(net4311),
    .B(_05319_),
    .Y(_05345_));
 NAND2x2_ASAP7_75t_R _11434_ (.A(net4311),
    .B(_05319_),
    .Y(_05346_));
 INVx1_ASAP7_75t_R _11435_ (.A(_05346_),
    .Y(_05347_));
 OAI21x1_ASAP7_75t_R _11436_ (.A1(_05345_),
    .A2(_05347_),
    .B(net2772),
    .Y(_05348_));
 INVx1_ASAP7_75t_R _11437_ (.A(_05348_),
    .Y(_05349_));
 NOR2x1_ASAP7_75t_R _11438_ (.A(net4613),
    .B(net4320),
    .Y(_05350_));
 XOR2x2_ASAP7_75t_R _11439_ (.A(_05350_),
    .B(net4671),
    .Y(_05351_));
 AND3x1_ASAP7_75t_R _11440_ (.A(_05351_),
    .B(_04436_),
    .C(net4936),
    .Y(_05352_));
 AND3x1_ASAP7_75t_R _11441_ (.A(_05344_),
    .B(_05349_),
    .C(_05352_),
    .Y(_05353_));
 AOI21x1_ASAP7_75t_R _11442_ (.A1(_05326_),
    .A2(_05353_),
    .B(net4320),
    .Y(_05354_));
 NAND2x2_ASAP7_75t_R _11443_ (.A(net5506),
    .B(_05354_),
    .Y(_05355_));
 BUFx3_ASAP7_75t_R place2950 (.A(_03967_),
    .Y(net2950));
 AOI21x1_ASAP7_75t_R _11445_ (.A1(net5591),
    .A2(_04335_),
    .B(net5359),
    .Y(_00808_));
 AO21x1_ASAP7_75t_R _11446_ (.A1(_05319_),
    .A2(net4256),
    .B(net2772),
    .Y(_05357_));
 AO21x1_ASAP7_75t_R _11447_ (.A1(_05339_),
    .A2(_05338_),
    .B(_05334_),
    .Y(_05358_));
 INVx1_ASAP7_75t_R _11448_ (.A(_05358_),
    .Y(_05359_));
 NAND2x1_ASAP7_75t_R _11449_ (.A(_05357_),
    .B(_05359_),
    .Y(_05360_));
 INVx1_ASAP7_75t_R _11450_ (.A(_05345_),
    .Y(_05361_));
 OA211x2_ASAP7_75t_R _11451_ (.A1(net4320),
    .A2(net4936),
    .B(net5019),
    .C(net4753),
    .Y(_05362_));
 OA21x2_ASAP7_75t_R _11452_ (.A1(net4362),
    .A2(net4670),
    .B(_05362_),
    .Y(_05363_));
 NAND2x1_ASAP7_75t_R _11453_ (.A(_05351_),
    .B(_05363_),
    .Y(_05364_));
 AO21x2_ASAP7_75t_R _11454_ (.A1(_05361_),
    .A2(net2734),
    .B(_05364_),
    .Y(_05365_));
 NOR2x1_ASAP7_75t_R _11455_ (.A(_05360_),
    .B(_05365_),
    .Y(_05366_));
 INVx1_ASAP7_75t_R _11456_ (.A(_05328_),
    .Y(_05367_));
 XOR2x2_ASAP7_75t_R _11457_ (.A(net2742),
    .B(_05367_),
    .Y(_05368_));
 NOR2x1_ASAP7_75t_R _11458_ (.A(_05368_),
    .B(_05325_),
    .Y(_05369_));
 AOI21x1_ASAP7_75t_R _11459_ (.A1(_05366_),
    .A2(_05369_),
    .B(net4320),
    .Y(_05370_));
 OAI21x1_ASAP7_75t_R _11460_ (.A1(net2706),
    .A2(net2699),
    .B(net5363),
    .Y(_05371_));
 AOI21x1_ASAP7_75t_R _11461_ (.A1(net5141),
    .A2(net5920),
    .B(_05371_),
    .Y(_00809_));
 NAND2x1p5_ASAP7_75t_R _11462_ (.A(net2700),
    .B(net4946),
    .Y(_05372_));
 BUFx3_ASAP7_75t_R place2949 (.A(_03967_),
    .Y(net2949));
 AOI21x1_ASAP7_75t_R _11464_ (.A1(net5591),
    .A2(_05372_),
    .B(net5359),
    .Y(_00810_));
 NAND2x2_ASAP7_75t_R _11465_ (.A(_05370_),
    .B(net5506),
    .Y(_05374_));
 NAND2x1p5_ASAP7_75t_R _11466_ (.A(net4947),
    .B(net2700),
    .Y(_05375_));
 AOI21x1_ASAP7_75t_R _11467_ (.A1(net2697),
    .A2(_05375_),
    .B(net5359),
    .Y(_00811_));
 BUFx3_ASAP7_75t_R place2946 (.A(_04021_),
    .Y(net2946));
 NAND2x1_ASAP7_75t_R _11469_ (.A(net5434),
    .B(net2700),
    .Y(_05377_));
 AOI21x1_ASAP7_75t_R _11470_ (.A1(net5591),
    .A2(_05377_),
    .B(net5359),
    .Y(_00812_));
 NAND2x1p5_ASAP7_75t_R _11471_ (.A(net4948),
    .B(net5920),
    .Y(_05378_));
 AOI21x1_ASAP7_75t_R _11472_ (.A1(net2697),
    .A2(_05378_),
    .B(net5359),
    .Y(_00813_));
 NAND2x1p5_ASAP7_75t_R _11473_ (.A(net4949),
    .B(net5920),
    .Y(_05379_));
 AOI21x1_ASAP7_75t_R _11474_ (.A1(net5591),
    .A2(_05379_),
    .B(net5359),
    .Y(_00814_));
 NAND2x1p5_ASAP7_75t_R _11475_ (.A(net4950),
    .B(net2700),
    .Y(_05380_));
 AOI21x1_ASAP7_75t_R _11476_ (.A1(net2697),
    .A2(_05380_),
    .B(net5359),
    .Y(_00815_));
 NAND2x1p5_ASAP7_75t_R _11477_ (.A(net4951),
    .B(net5920),
    .Y(_05381_));
 AOI21x1_ASAP7_75t_R _11478_ (.A1(net5591),
    .A2(_05381_),
    .B(net5359),
    .Y(_00816_));
 NAND2x1p5_ASAP7_75t_R _11479_ (.A(net4952),
    .B(net2700),
    .Y(_05382_));
 AOI21x1_ASAP7_75t_R _11480_ (.A1(net2698),
    .A2(_05382_),
    .B(net5359),
    .Y(_00817_));
 AO21x1_ASAP7_75t_R _11481_ (.A1(net4753),
    .A2(net2710),
    .B(net5359),
    .Y(_05383_));
 AOI21x1_ASAP7_75t_R _11482_ (.A1(net5132),
    .A2(net5923),
    .B(_05383_),
    .Y(_00818_));
 NAND2x1p5_ASAP7_75t_R _11483_ (.A(net4953),
    .B(net2701),
    .Y(_05384_));
 AOI21x1_ASAP7_75t_R _11484_ (.A1(net2696),
    .A2(_05384_),
    .B(net5359),
    .Y(_00819_));
 NAND2x1p5_ASAP7_75t_R _11485_ (.A(net4954),
    .B(net5912),
    .Y(_05385_));
 AOI21x1_ASAP7_75t_R _11486_ (.A1(net2698),
    .A2(_05385_),
    .B(net5359),
    .Y(_00820_));
 NAND2x1p5_ASAP7_75t_R _11487_ (.A(net5912),
    .B(net4955),
    .Y(_05386_));
 BUFx3_ASAP7_75t_R place2944 (.A(_05200_),
    .Y(net2944));
 AOI21x1_ASAP7_75t_R _11489_ (.A1(net2696),
    .A2(_05386_),
    .B(net5359),
    .Y(_00821_));
 NAND2x1p5_ASAP7_75t_R _11490_ (.A(net2702),
    .B(net4956),
    .Y(_05388_));
 AOI21x1_ASAP7_75t_R _11491_ (.A1(net2698),
    .A2(_05388_),
    .B(net5359),
    .Y(_00822_));
 NAND2x1p5_ASAP7_75t_R _11492_ (.A(net5912),
    .B(net4957),
    .Y(_05389_));
 AOI21x1_ASAP7_75t_R _11493_ (.A1(net2696),
    .A2(_05389_),
    .B(net5359),
    .Y(_00823_));
 NAND2x1p5_ASAP7_75t_R _11494_ (.A(net2702),
    .B(net4958),
    .Y(_05390_));
 AOI21x1_ASAP7_75t_R _11495_ (.A1(net2698),
    .A2(_05390_),
    .B(net5359),
    .Y(_00824_));
 NAND2x1p5_ASAP7_75t_R _11496_ (.A(net2702),
    .B(net4959),
    .Y(_05391_));
 AOI21x1_ASAP7_75t_R _11497_ (.A1(net2696),
    .A2(_05391_),
    .B(net5359),
    .Y(_00825_));
 NAND2x1p5_ASAP7_75t_R _11498_ (.A(net4960),
    .B(net2702),
    .Y(_05392_));
 AOI21x1_ASAP7_75t_R _11499_ (.A1(net2698),
    .A2(_05392_),
    .B(net5359),
    .Y(_00826_));
 NAND2x1p5_ASAP7_75t_R _11500_ (.A(net5912),
    .B(net4961),
    .Y(_05393_));
 AOI21x1_ASAP7_75t_R _11501_ (.A1(net2696),
    .A2(_05393_),
    .B(net5359),
    .Y(_00827_));
 NAND2x1p5_ASAP7_75t_R _11502_ (.A(net4962),
    .B(net2702),
    .Y(_05394_));
 AOI21x1_ASAP7_75t_R _11503_ (.A1(net2698),
    .A2(_05394_),
    .B(net5359),
    .Y(_00828_));
 AO21x1_ASAP7_75t_R _11504_ (.A1(net4670),
    .A2(net2710),
    .B(net5359),
    .Y(_05395_));
 AOI21x1_ASAP7_75t_R _11505_ (.A1(net5923),
    .A2(net5124),
    .B(_05395_),
    .Y(_00829_));
 NAND2x1p5_ASAP7_75t_R _11506_ (.A(net4963),
    .B(net5912),
    .Y(_05396_));
 AOI21x1_ASAP7_75t_R _11507_ (.A1(net2696),
    .A2(_05396_),
    .B(net5359),
    .Y(_00830_));
 NAND2x1p5_ASAP7_75t_R _11508_ (.A(net4882),
    .B(net2700),
    .Y(_05397_));
 AOI21x1_ASAP7_75t_R _11509_ (.A1(net2697),
    .A2(_05397_),
    .B(net5359),
    .Y(_00831_));
 NOR2x1_ASAP7_75t_R _11510_ (.A(net4320),
    .B(_05363_),
    .Y(_05398_));
 XOR2x2_ASAP7_75t_R _11511_ (.A(_05398_),
    .B(net4191),
    .Y(_05399_));
 NOR2x1p5_ASAP7_75t_R _11512_ (.A(net4937),
    .B(net2710),
    .Y(_05400_));
 AOI211x1_ASAP7_75t_R _11513_ (.A1(net2710),
    .A2(_05399_),
    .B(_05400_),
    .C(net5359),
    .Y(_00832_));
 NAND2x1_ASAP7_75t_R _11514_ (.A(net2735),
    .B(net2729),
    .Y(_05401_));
 NOR2x1_ASAP7_75t_R _11515_ (.A(net4320),
    .B(_05352_),
    .Y(_05402_));
 XOR2x2_ASAP7_75t_R _11516_ (.A(_05401_),
    .B(_05402_),
    .Y(_05403_));
 NOR2x1p5_ASAP7_75t_R _11517_ (.A(net4938),
    .B(net5540),
    .Y(_05404_));
 AOI211x1_ASAP7_75t_R _11518_ (.A1(net5540),
    .A2(_05403_),
    .B(_05404_),
    .C(net5359),
    .Y(_00833_));
 AND2x2_ASAP7_75t_R _11519_ (.A(_05357_),
    .B(net2736),
    .Y(_05405_));
 NAND2x1_ASAP7_75t_R _11520_ (.A(net4362),
    .B(net2719),
    .Y(_05406_));
 XNOR2x2_ASAP7_75t_R _11521_ (.A(_05405_),
    .B(_05406_),
    .Y(_05407_));
 AO21x1_ASAP7_75t_R _11522_ (.A1(_05407_),
    .A2(net5541),
    .B(net5359),
    .Y(_05408_));
 AOI21x1_ASAP7_75t_R _11523_ (.A1(net5121),
    .A2(net2699),
    .B(_05408_),
    .Y(_00834_));
 AO21x1_ASAP7_75t_R _11524_ (.A1(_05349_),
    .A2(_05352_),
    .B(net4320),
    .Y(_05409_));
 XNOR2x2_ASAP7_75t_R _11525_ (.A(net2730),
    .B(_05409_),
    .Y(_05410_));
 NOR2x1p5_ASAP7_75t_R _11526_ (.A(net4940),
    .B(net5538),
    .Y(_05411_));
 AOI211x1_ASAP7_75t_R _11527_ (.A1(_05410_),
    .A2(net5538),
    .B(_05411_),
    .C(net5359),
    .Y(_00835_));
 OAI21x1_ASAP7_75t_R _11528_ (.A1(net2720),
    .A2(net2719),
    .B(net4362),
    .Y(_05412_));
 XOR2x2_ASAP7_75t_R _11529_ (.A(_05412_),
    .B(net2737),
    .Y(_05413_));
 OAI21x1_ASAP7_75t_R _11530_ (.A1(net2699),
    .A2(_05413_),
    .B(net5363),
    .Y(_05414_));
 AOI21x1_ASAP7_75t_R _11531_ (.A1(net5119),
    .A2(net5920),
    .B(_05414_),
    .Y(_00836_));
 NAND2x1p5_ASAP7_75t_R _11532_ (.A(net4942),
    .B(net5920),
    .Y(_05415_));
 INVx1_ASAP7_75t_R _11533_ (.A(_05402_),
    .Y(_05416_));
 OAI21x1_ASAP7_75t_R _11534_ (.A1(net2721),
    .A2(net2722),
    .B(net4362),
    .Y(_05417_));
 AOI21x1_ASAP7_75t_R _11535_ (.A1(_05416_),
    .A2(_05417_),
    .B(net2731),
    .Y(_05418_));
 AND3x1_ASAP7_75t_R _11536_ (.A(_05417_),
    .B(net2731),
    .C(_05416_),
    .Y(_05419_));
 OAI21x1_ASAP7_75t_R _11537_ (.A1(_05418_),
    .A2(_05419_),
    .B(net5539),
    .Y(_05420_));
 AOI21x1_ASAP7_75t_R _11538_ (.A1(_05420_),
    .A2(_05415_),
    .B(net5359),
    .Y(_00837_));
 AOI21x1_ASAP7_75t_R _11539_ (.A1(net5117),
    .A2(net5920),
    .B(_05371_),
    .Y(_00838_));
 NOR2x1_ASAP7_75t_R _11540_ (.A(net5360),
    .B(net5033),
    .Y(_00839_));
 NAND2x1_ASAP7_75t_R _11541_ (.A(net5024),
    .B(net5021),
    .Y(_05421_));
 NAND2x1p5_ASAP7_75t_R _11542_ (.A(net5200),
    .B(net5635),
    .Y(_05422_));
 AND3x1_ASAP7_75t_R _11543_ (.A(_05422_),
    .B(net5363),
    .C(_05421_),
    .Y(_00840_));
 BUFx3_ASAP7_75t_R place2942 (.A(_05202_),
    .Y(net2942));
 OR3x1_ASAP7_75t_R _11545_ (.A(_00070_),
    .B(_00060_),
    .C(_00541_),
    .Y(_05424_));
 NOR3x1_ASAP7_75t_R _11546_ (.A(_05424_),
    .B(_00025_),
    .C(_00026_),
    .Y(_05425_));
 INVx1_ASAP7_75t_R _11547_ (.A(_00027_),
    .Y(_05426_));
 INVx1_ASAP7_75t_R _11548_ (.A(_00028_),
    .Y(_05427_));
 AND3x4_ASAP7_75t_R _11549_ (.A(_05426_),
    .B(_05425_),
    .C(_05427_),
    .Y(_05428_));
 XOR2x2_ASAP7_75t_R _11550_ (.A(net4607),
    .B(net5013),
    .Y(_05429_));
 INVx1_ASAP7_75t_R _11551_ (.A(_05429_),
    .Y(_05430_));
 OR3x1_ASAP7_75t_R _11552_ (.A(_00060_),
    .B(net5115),
    .C(net5104),
    .Y(_05431_));
 XOR2x2_ASAP7_75t_R _11553_ (.A(_05431_),
    .B(net5089),
    .Y(_05432_));
 INVx2_ASAP7_75t_R _11554_ (.A(_05432_),
    .Y(_05433_));
 XOR2x2_ASAP7_75t_R _11555_ (.A(net4722),
    .B(net5088),
    .Y(_05434_));
 INVx1_ASAP7_75t_R _11556_ (.A(_05434_),
    .Y(_05435_));
 XOR2x2_ASAP7_75t_R _11557_ (.A(net4815),
    .B(net5093),
    .Y(_05436_));
 INVx1_ASAP7_75t_R _11558_ (.A(_05436_),
    .Y(_05437_));
 AND3x1_ASAP7_75t_R _11559_ (.A(_05437_),
    .B(_00542_),
    .C(net5021),
    .Y(_05438_));
 AND3x1_ASAP7_75t_R _11560_ (.A(net4721),
    .B(net4606),
    .C(_05438_),
    .Y(_05439_));
 NOR3x1_ASAP7_75t_R _11561_ (.A(_05431_),
    .B(_00025_),
    .C(net5089),
    .Y(_05440_));
 XOR2x2_ASAP7_75t_R _11562_ (.A(_05440_),
    .B(_02426_),
    .Y(_05441_));
 INVx1_ASAP7_75t_R _11563_ (.A(_05441_),
    .Y(_05442_));
 XOR2x2_ASAP7_75t_R _11564_ (.A(net4666),
    .B(net5086),
    .Y(_05443_));
 AND3x1_ASAP7_75t_R _11565_ (.A(_05439_),
    .B(net4663),
    .C(net4605),
    .Y(_05444_));
 AND3x4_ASAP7_75t_R _11566_ (.A(_05426_),
    .B(_02426_),
    .C(_05440_),
    .Y(_05445_));
 XOR2x2_ASAP7_75t_R _11567_ (.A(_05445_),
    .B(_05427_),
    .Y(_05446_));
 INVx1_ASAP7_75t_R _11568_ (.A(_05446_),
    .Y(_05447_));
 AND2x2_ASAP7_75t_R _11569_ (.A(_05444_),
    .B(net4604),
    .Y(_05448_));
 INVx1_ASAP7_75t_R _11570_ (.A(_00053_),
    .Y(_05449_));
 INVx1_ASAP7_75t_R _11571_ (.A(net5100),
    .Y(_05450_));
 NOR2x1_ASAP7_75t_R _11572_ (.A(_00031_),
    .B(_00030_),
    .Y(_05451_));
 AND3x1_ASAP7_75t_R _11573_ (.A(net4878),
    .B(_05427_),
    .C(net5013),
    .Y(_05452_));
 INVx1_ASAP7_75t_R _11574_ (.A(_00033_),
    .Y(_05453_));
 INVx1_ASAP7_75t_R _11575_ (.A(_00035_),
    .Y(_05454_));
 AND5x2_ASAP7_75t_R _11576_ (.A(_05452_),
    .B(net5015),
    .C(net4877),
    .D(net5009),
    .E(net4876),
    .Y(_05455_));
 INVx1_ASAP7_75t_R _11577_ (.A(_00038_),
    .Y(_05456_));
 INVx1_ASAP7_75t_R _11578_ (.A(_00039_),
    .Y(_05457_));
 AND4x1_ASAP7_75t_R _11579_ (.A(net5010),
    .B(_02477_),
    .C(_05456_),
    .D(_05457_),
    .Y(_05458_));
 NOR2x1_ASAP7_75t_R _11580_ (.A(_00040_),
    .B(_00041_),
    .Y(_05459_));
 INVx1_ASAP7_75t_R _11581_ (.A(_00042_),
    .Y(_05460_));
 AND3x1_ASAP7_75t_R _11582_ (.A(_05459_),
    .B(_05460_),
    .C(_02487_),
    .Y(_05461_));
 AND2x2_ASAP7_75t_R _11583_ (.A(_05458_),
    .B(_05461_),
    .Y(_05462_));
 AND5x2_ASAP7_75t_R _11584_ (.A(net4719),
    .B(_05455_),
    .C(_05462_),
    .D(_02458_),
    .E(_05450_),
    .Y(_05463_));
 INVx1_ASAP7_75t_R _11585_ (.A(net5097),
    .Y(_05464_));
 AND3x4_ASAP7_75t_R _11586_ (.A(_02454_),
    .B(_05464_),
    .C(_05463_),
    .Y(_05465_));
 INVx1_ASAP7_75t_R _11587_ (.A(_00051_),
    .Y(_05466_));
 NOR2x1_ASAP7_75t_R _11588_ (.A(net5095),
    .B(_00050_),
    .Y(_05467_));
 AND4x2_ASAP7_75t_R _11589_ (.A(_05465_),
    .B(_05466_),
    .C(_02463_),
    .D(_05467_),
    .Y(_05468_));
 NOR2x1p5_ASAP7_75t_R _11590_ (.A(_05449_),
    .B(_05468_),
    .Y(_05469_));
 AND2x4_ASAP7_75t_R _11591_ (.A(_05468_),
    .B(_05449_),
    .Y(_05470_));
 NOR2x2_ASAP7_75t_R _11592_ (.A(_05469_),
    .B(_05470_),
    .Y(_05471_));
 INVx3_ASAP7_75t_R _11593_ (.A(_05471_),
    .Y(_05472_));
 BUFx3_ASAP7_75t_R place2941 (.A(_05245_),
    .Y(net2941));
 AO21x1_ASAP7_75t_R _11595_ (.A1(net4508),
    .A2(_05448_),
    .B(net4400),
    .Y(_05474_));
 AND3x1_ASAP7_75t_R _11596_ (.A(_05445_),
    .B(_05427_),
    .C(net5013),
    .Y(_05475_));
 XOR2x2_ASAP7_75t_R _11597_ (.A(_05475_),
    .B(_02392_),
    .Y(_05476_));
 XOR2x2_ASAP7_75t_R _11598_ (.A(_05474_),
    .B(net4603),
    .Y(_05477_));
 INVx1_ASAP7_75t_R _11599_ (.A(_05477_),
    .Y(_05478_));
 NOR2x1_ASAP7_75t_R _11600_ (.A(_05429_),
    .B(_05476_),
    .Y(_05479_));
 INVx1_ASAP7_75t_R _11601_ (.A(net5093),
    .Y(_05480_));
 INVx1_ASAP7_75t_R _11602_ (.A(net4815),
    .Y(_05481_));
 AND3x1_ASAP7_75t_R _11603_ (.A(_05433_),
    .B(_05480_),
    .C(_05481_),
    .Y(_05482_));
 AND3x1_ASAP7_75t_R _11604_ (.A(_05442_),
    .B(_05482_),
    .C(_05435_),
    .Y(_05483_));
 AND3x1_ASAP7_75t_R _11605_ (.A(_05443_),
    .B(_05483_),
    .C(_05447_),
    .Y(_05484_));
 AND2x2_ASAP7_75t_R _11606_ (.A(_05484_),
    .B(_05479_),
    .Y(_05485_));
 NOR2x1_ASAP7_75t_R _11607_ (.A(net4454),
    .B(net4400),
    .Y(_05486_));
 NAND3x1_ASAP7_75t_R _11608_ (.A(net4607),
    .B(net5013),
    .C(_02392_),
    .Y(_05487_));
 XOR2x2_ASAP7_75t_R _11609_ (.A(_05487_),
    .B(net5114),
    .Y(_05488_));
 INVx1_ASAP7_75t_R _11610_ (.A(_05488_),
    .Y(_05489_));
 XOR2x2_ASAP7_75t_R _11611_ (.A(_05486_),
    .B(net4453),
    .Y(_05490_));
 INVx1_ASAP7_75t_R _11612_ (.A(_05490_),
    .Y(_05491_));
 AND3x1_ASAP7_75t_R _11613_ (.A(_05455_),
    .B(net4719),
    .C(_05458_),
    .Y(_05492_));
 AND2x2_ASAP7_75t_R _11614_ (.A(_05492_),
    .B(net4874),
    .Y(_05493_));
 XOR2x2_ASAP7_75t_R _11615_ (.A(_05493_),
    .B(net4873),
    .Y(_05494_));
 AND3x1_ASAP7_75t_R _11616_ (.A(_05451_),
    .B(_02407_),
    .C(_02389_),
    .Y(_05495_));
 AND3x1_ASAP7_75t_R _11617_ (.A(_05495_),
    .B(_05453_),
    .C(_02449_),
    .Y(_05496_));
 AND3x1_ASAP7_75t_R _11618_ (.A(_05496_),
    .B(_05454_),
    .C(_02445_),
    .Y(_05497_));
 NAND2x1p5_ASAP7_75t_R _11619_ (.A(_05428_),
    .B(_05497_),
    .Y(_05498_));
 OR3x1_ASAP7_75t_R _11620_ (.A(net5108),
    .B(_05498_),
    .C(net5107),
    .Y(_05499_));
 OR3x1_ASAP7_75t_R _11621_ (.A(net5106),
    .B(_05499_),
    .C(net5105),
    .Y(_05500_));
 OR3x1_ASAP7_75t_R _11622_ (.A(net5102),
    .B(net5103),
    .C(_05500_),
    .Y(_05501_));
 XOR2x2_ASAP7_75t_R _11623_ (.A(net5101),
    .B(_05501_),
    .Y(_05502_));
 NOR2x1p5_ASAP7_75t_R _11624_ (.A(_05494_),
    .B(_05502_),
    .Y(_05503_));
 XOR2x2_ASAP7_75t_R _11625_ (.A(net4500),
    .B(net5106),
    .Y(_05504_));
 INVx1_ASAP7_75t_R _11626_ (.A(_05504_),
    .Y(_05505_));
 XOR2x2_ASAP7_75t_R _11627_ (.A(net4545),
    .B(net5108),
    .Y(_05506_));
 NAND2x1_ASAP7_75t_R _11628_ (.A(net4719),
    .B(_05455_),
    .Y(_05507_));
 XOR2x2_ASAP7_75t_R _11629_ (.A(net4660),
    .B(net5109),
    .Y(_05508_));
 NOR2x1_ASAP7_75t_R _11630_ (.A(_05506_),
    .B(_05508_),
    .Y(_05509_));
 OR3x1_ASAP7_75t_R _11631_ (.A(_05507_),
    .B(net5109),
    .C(net5108),
    .Y(_05510_));
 XOR2x2_ASAP7_75t_R _11632_ (.A(_05510_),
    .B(net4875),
    .Y(_05511_));
 AND3x1_ASAP7_75t_R _11633_ (.A(_05505_),
    .B(_05509_),
    .C(_05511_),
    .Y(_05512_));
 XNOR2x2_ASAP7_75t_R _11634_ (.A(net5105),
    .B(_05492_),
    .Y(_05513_));
 XOR2x2_ASAP7_75t_R _11635_ (.A(_05500_),
    .B(net5103),
    .Y(_05514_));
 NOR2x1_ASAP7_75t_R _11636_ (.A(_05513_),
    .B(_05514_),
    .Y(_05515_));
 AND3x1_ASAP7_75t_R _11637_ (.A(net4306),
    .B(net4348),
    .C(_05515_),
    .Y(_05516_));
 INVx1_ASAP7_75t_R _11638_ (.A(_05516_),
    .Y(_05517_));
 OR4x1_ASAP7_75t_R _11639_ (.A(net5103),
    .B(net5102),
    .C(net5101),
    .D(_00044_),
    .Y(_05518_));
 OR4x1_ASAP7_75t_R _11640_ (.A(_05499_),
    .B(net5106),
    .C(net5105),
    .D(_05518_),
    .Y(_05519_));
 NOR2x1_ASAP7_75t_R _11641_ (.A(net5099),
    .B(net4450),
    .Y(_05520_));
 AO21x1_ASAP7_75t_R _11642_ (.A1(_05520_),
    .A2(net4872),
    .B(net5008),
    .Y(_05521_));
 OR4x1_ASAP7_75t_R _11643_ (.A(_05519_),
    .B(net5099),
    .C(net5098),
    .D(net5096),
    .Y(_05522_));
 NAND2x1_ASAP7_75t_R _11644_ (.A(_05521_),
    .B(_05522_),
    .Y(_05523_));
 NOR2x1_ASAP7_75t_R _11645_ (.A(net4872),
    .B(net4662),
    .Y(_05524_));
 AND2x2_ASAP7_75t_R _11646_ (.A(net4662),
    .B(net4872),
    .Y(_05525_));
 NOR2x1_ASAP7_75t_R _11647_ (.A(_05524_),
    .B(_05525_),
    .Y(_05526_));
 INVx1_ASAP7_75t_R _11648_ (.A(_05526_),
    .Y(_05527_));
 NAND2x1_ASAP7_75t_R _11649_ (.A(_05461_),
    .B(_05492_),
    .Y(_05528_));
 XOR2x2_ASAP7_75t_R _11650_ (.A(_05528_),
    .B(net5100),
    .Y(_05529_));
 XOR2x2_ASAP7_75t_R _11651_ (.A(net4450),
    .B(net5099),
    .Y(_05530_));
 NOR2x1_ASAP7_75t_R _11652_ (.A(_05529_),
    .B(_05530_),
    .Y(_05531_));
 AND3x1_ASAP7_75t_R _11653_ (.A(_05523_),
    .B(_05527_),
    .C(_05531_),
    .Y(_05532_));
 XNOR2x2_ASAP7_75t_R _11654_ (.A(net5095),
    .B(_05465_),
    .Y(_05533_));
 OR5x1_ASAP7_75t_R _11655_ (.A(net5099),
    .B(_05518_),
    .C(_00047_),
    .D(_00048_),
    .E(_00049_),
    .Y(_05534_));
 NOR2x1_ASAP7_75t_R _11656_ (.A(_05534_),
    .B(_05500_),
    .Y(_05535_));
 NOR2x1_ASAP7_75t_R _11657_ (.A(_02469_),
    .B(net4395),
    .Y(_05536_));
 INVx1_ASAP7_75t_R _11658_ (.A(_05536_),
    .Y(_05537_));
 AND2x2_ASAP7_75t_R _11659_ (.A(_05535_),
    .B(_02469_),
    .Y(_05538_));
 INVx1_ASAP7_75t_R _11660_ (.A(_05538_),
    .Y(_05539_));
 NAND2x1p5_ASAP7_75t_R _11661_ (.A(_05537_),
    .B(_05539_),
    .Y(_05540_));
 INVx1_ASAP7_75t_R _11662_ (.A(_05540_),
    .Y(_05541_));
 NOR2x1_ASAP7_75t_R _11663_ (.A(_05533_),
    .B(_05541_),
    .Y(_05542_));
 INVx1_ASAP7_75t_R _11664_ (.A(_05542_),
    .Y(_05543_));
 NAND2x1_ASAP7_75t_R _11665_ (.A(net4872),
    .B(_05520_),
    .Y(_05544_));
 NAND2x1_ASAP7_75t_R _11666_ (.A(_05466_),
    .B(_05467_),
    .Y(_05545_));
 NOR3x1_ASAP7_75t_R _11667_ (.A(_05544_),
    .B(net5096),
    .C(_05545_),
    .Y(_05546_));
 NOR2x1_ASAP7_75t_R _11668_ (.A(net5006),
    .B(_05546_),
    .Y(_05547_));
 INVx1_ASAP7_75t_R _11669_ (.A(_05546_),
    .Y(_05548_));
 NOR2x1_ASAP7_75t_R _11670_ (.A(net5091),
    .B(_05548_),
    .Y(_05549_));
 AND4x1_ASAP7_75t_R _11671_ (.A(net4662),
    .B(net4872),
    .C(net5008),
    .D(_05467_),
    .Y(_05550_));
 XOR2x2_ASAP7_75t_R _11672_ (.A(_05550_),
    .B(net5094),
    .Y(_05551_));
 OAI21x1_ASAP7_75t_R _11673_ (.A1(_05547_),
    .A2(_05549_),
    .B(net4540),
    .Y(_05552_));
 NOR2x1_ASAP7_75t_R _11674_ (.A(_05543_),
    .B(_05552_),
    .Y(_05553_));
 NAND2x1_ASAP7_75t_R _11675_ (.A(_05532_),
    .B(_05553_),
    .Y(_05554_));
 NOR2x1_ASAP7_75t_R _11676_ (.A(_05517_),
    .B(_05554_),
    .Y(_05555_));
 AND2x2_ASAP7_75t_R _11677_ (.A(net4607),
    .B(net4718),
    .Y(_05556_));
 XOR2x2_ASAP7_75t_R _11678_ (.A(_05556_),
    .B(net4876),
    .Y(_05557_));
 AND2x2_ASAP7_75t_R _11679_ (.A(_05475_),
    .B(net4878),
    .Y(_05558_));
 INVx1_ASAP7_75t_R _11680_ (.A(_05558_),
    .Y(_05559_));
 OR3x1_ASAP7_75t_R _11681_ (.A(_05559_),
    .B(net5113),
    .C(net5112),
    .Y(_05560_));
 XOR2x2_ASAP7_75t_R _11682_ (.A(_05560_),
    .B(net5111),
    .Y(_05561_));
 NOR2x1_ASAP7_75t_R _11683_ (.A(_05557_),
    .B(net4449),
    .Y(_05562_));
 NOR2x1_ASAP7_75t_R _11684_ (.A(net4501),
    .B(net4603),
    .Y(_05563_));
 AND3x1_ASAP7_75t_R _11685_ (.A(_05563_),
    .B(_05430_),
    .C(net4604),
    .Y(_05564_));
 XOR2x2_ASAP7_75t_R _11686_ (.A(net4600),
    .B(net5113),
    .Y(_05565_));
 AND2x2_ASAP7_75t_R _11687_ (.A(net4607),
    .B(net4836),
    .Y(_05566_));
 XOR2x2_ASAP7_75t_R _11688_ (.A(_05566_),
    .B(net5112),
    .Y(_05567_));
 AND2x2_ASAP7_75t_R _11689_ (.A(net4539),
    .B(_05567_),
    .Y(_05568_));
 AND4x1_ASAP7_75t_R _11690_ (.A(net4394),
    .B(net4507),
    .C(net4393),
    .D(_05568_),
    .Y(_05569_));
 NAND3x1_ASAP7_75t_R _11691_ (.A(net4455),
    .B(_05555_),
    .C(_05569_),
    .Y(_05570_));
 INVx1_ASAP7_75t_R _11692_ (.A(_05570_),
    .Y(_05571_));
 NOR2x1_ASAP7_75t_R _11693_ (.A(net4251),
    .B(net4190),
    .Y(_05572_));
 INVx1_ASAP7_75t_R _11694_ (.A(_05572_),
    .Y(_05573_));
 AND3x1_ASAP7_75t_R _11695_ (.A(_05485_),
    .B(_05565_),
    .C(_05489_),
    .Y(_05574_));
 INVx1_ASAP7_75t_R _11696_ (.A(_05561_),
    .Y(_05575_));
 AND3x2_ASAP7_75t_R _11697_ (.A(_05574_),
    .B(_05575_),
    .C(_05567_),
    .Y(_05576_));
 INVx1_ASAP7_75t_R _11698_ (.A(_05523_),
    .Y(_05577_));
 NAND2x1_ASAP7_75t_R _11699_ (.A(_05540_),
    .B(_05551_),
    .Y(_05578_));
 NOR3x1_ASAP7_75t_R _11700_ (.A(_05577_),
    .B(_05533_),
    .C(_05578_),
    .Y(_05579_));
 NOR2x1_ASAP7_75t_R _11701_ (.A(_05494_),
    .B(_05514_),
    .Y(_05580_));
 NOR2x1_ASAP7_75t_R _11702_ (.A(_05513_),
    .B(net4452),
    .Y(_05581_));
 INVx1_ASAP7_75t_R _11703_ (.A(_05511_),
    .Y(_05582_));
 NOR2x1_ASAP7_75t_R _11704_ (.A(net4498),
    .B(_05582_),
    .Y(_05583_));
 NOR2x1_ASAP7_75t_R _11705_ (.A(_05557_),
    .B(_05508_),
    .Y(_05584_));
 AND2x2_ASAP7_75t_R _11706_ (.A(_05583_),
    .B(_05584_),
    .Y(_05585_));
 AND3x1_ASAP7_75t_R _11707_ (.A(_05580_),
    .B(_05581_),
    .C(_05585_),
    .Y(_05586_));
 NOR2x1_ASAP7_75t_R _11708_ (.A(net4543),
    .B(_05502_),
    .Y(_05587_));
 NOR2x1_ASAP7_75t_R _11709_ (.A(net4544),
    .B(net4396),
    .Y(_05588_));
 AND2x2_ASAP7_75t_R _11710_ (.A(_05587_),
    .B(_05588_),
    .Y(_05589_));
 AND3x1_ASAP7_75t_R _11711_ (.A(_05579_),
    .B(_05586_),
    .C(_05589_),
    .Y(_05590_));
 AOI21x1_ASAP7_75t_R _11712_ (.A1(net4345),
    .A2(_05590_),
    .B(_05472_),
    .Y(_05591_));
 NOR2x1_ASAP7_75t_R _11713_ (.A(_05573_),
    .B(_05591_),
    .Y(_05592_));
 NAND2x1_ASAP7_75t_R _11714_ (.A(_05573_),
    .B(_05591_),
    .Y(_05593_));
 INVx1_ASAP7_75t_R _11715_ (.A(_05593_),
    .Y(_05594_));
 NOR2x1_ASAP7_75t_R _11716_ (.A(net4005),
    .B(_05594_),
    .Y(_05595_));
 NOR2x1_ASAP7_75t_R _11717_ (.A(_05571_),
    .B(_05595_),
    .Y(_05596_));
 INVx1_ASAP7_75t_R _11718_ (.A(_05596_),
    .Y(_05597_));
 OR3x1_ASAP7_75t_R _11719_ (.A(net4504),
    .B(net4505),
    .C(_05588_),
    .Y(_05598_));
 AND3x2_ASAP7_75t_R _11720_ (.A(_05576_),
    .B(_05583_),
    .C(_05584_),
    .Y(_05599_));
 AND2x2_ASAP7_75t_R _11721_ (.A(_05580_),
    .B(_05581_),
    .Y(_05600_));
 AND2x2_ASAP7_75t_R _11722_ (.A(_05599_),
    .B(_05600_),
    .Y(_05601_));
 AO21x1_ASAP7_75t_R _11723_ (.A1(_05601_),
    .A2(_05587_),
    .B(_05472_),
    .Y(_05602_));
 NAND2x1_ASAP7_75t_R _11724_ (.A(net4304),
    .B(net4188),
    .Y(_05603_));
 XOR2x2_ASAP7_75t_R _11725_ (.A(_05603_),
    .B(net4250),
    .Y(_05604_));
 INVx1_ASAP7_75t_R _11726_ (.A(_05592_),
    .Y(_05605_));
 AOI21x1_ASAP7_75t_R _11727_ (.A1(_05593_),
    .A2(_05605_),
    .B(_05570_),
    .Y(_05606_));
 INVx1_ASAP7_75t_R _11728_ (.A(_05606_),
    .Y(_05607_));
 AND2x2_ASAP7_75t_R _11729_ (.A(net4663),
    .B(net4605),
    .Y(_05608_));
 AND5x1_ASAP7_75t_R _11730_ (.A(net4721),
    .B(_05564_),
    .C(_05438_),
    .D(net4606),
    .E(_05608_),
    .Y(_05609_));
 AND3x1_ASAP7_75t_R _11731_ (.A(_05562_),
    .B(_05568_),
    .C(_05512_),
    .Y(_05610_));
 AND2x2_ASAP7_75t_R _11732_ (.A(_05503_),
    .B(_05515_),
    .Y(_05611_));
 AND3x1_ASAP7_75t_R _11733_ (.A(_05532_),
    .B(_05610_),
    .C(_05611_),
    .Y(_05612_));
 NAND2x1p5_ASAP7_75t_R _11734_ (.A(_05609_),
    .B(_05612_),
    .Y(_05613_));
 XOR2x2_ASAP7_75t_R _11735_ (.A(_05613_),
    .B(net4542),
    .Y(_05614_));
 INVx1_ASAP7_75t_R _11736_ (.A(net4542),
    .Y(_05615_));
 NAND2x1_ASAP7_75t_R _11737_ (.A(net4495),
    .B(net4401),
    .Y(_05616_));
 OAI21x1_ASAP7_75t_R _11738_ (.A1(net4401),
    .A2(_05614_),
    .B(_05616_),
    .Y(_05617_));
 AO21x1_ASAP7_75t_R _11739_ (.A1(net4305),
    .A2(_05615_),
    .B(_05472_),
    .Y(_05618_));
 NAND3x1_ASAP7_75t_R _11740_ (.A(_05602_),
    .B(_05598_),
    .C(_05618_),
    .Y(_05619_));
 XOR2x2_ASAP7_75t_R _11741_ (.A(net4252),
    .B(_05619_),
    .Y(_05620_));
 NAND3x1_ASAP7_75t_R _11742_ (.A(_05607_),
    .B(_05617_),
    .C(net5655),
    .Y(_05621_));
 AND5x1_ASAP7_75t_R _11743_ (.A(_05562_),
    .B(_05515_),
    .C(net4399),
    .D(net4451),
    .E(_05511_),
    .Y(_05622_));
 AND2x2_ASAP7_75t_R _11744_ (.A(net4306),
    .B(net4346),
    .Y(_05623_));
 AND3x1_ASAP7_75t_R _11745_ (.A(_05542_),
    .B(_05523_),
    .C(_05527_),
    .Y(_05624_));
 AND3x1_ASAP7_75t_R _11746_ (.A(_05430_),
    .B(net4604),
    .C(_05608_),
    .Y(_05625_));
 AND4x1_ASAP7_75t_R _11747_ (.A(_05568_),
    .B(net4548),
    .C(_05563_),
    .D(_05625_),
    .Y(_05626_));
 AND4x1_ASAP7_75t_R _11748_ (.A(_05622_),
    .B(_05623_),
    .C(_05624_),
    .D(_05626_),
    .Y(_05627_));
 XNOR2x2_ASAP7_75t_R _11749_ (.A(net4541),
    .B(_05627_),
    .Y(_05628_));
 BUFx3_ASAP7_75t_R place2940 (.A(_06288_),
    .Y(net2940));
 AND2x2_ASAP7_75t_R _11751_ (.A(net4401),
    .B(net4541),
    .Y(_05630_));
 AO21x2_ASAP7_75t_R _11752_ (.A1(_05628_),
    .A2(net4456),
    .B(_05630_),
    .Y(_05631_));
 INVx2_ASAP7_75t_R _11753_ (.A(_05631_),
    .Y(_05632_));
 OAI21x1_ASAP7_75t_R _11754_ (.A1(_05604_),
    .A2(_05621_),
    .B(_05632_),
    .Y(_05633_));
 AND2x2_ASAP7_75t_R _11755_ (.A(_05595_),
    .B(_05571_),
    .Y(_05634_));
 INVx1_ASAP7_75t_R _11756_ (.A(_05634_),
    .Y(_05635_));
 OAI21x1_ASAP7_75t_R _11757_ (.A1(_05633_),
    .A2(_05597_),
    .B(_05635_),
    .Y(_05636_));
 INVx2_ASAP7_75t_R _11758_ (.A(_05604_),
    .Y(_05637_));
 NAND2x1_ASAP7_75t_R _11759_ (.A(net4032),
    .B(net3967),
    .Y(_05638_));
 INVx1_ASAP7_75t_R _11760_ (.A(net3956),
    .Y(_05639_));
 AND3x1_ASAP7_75t_R _11761_ (.A(net3938),
    .B(net4031),
    .C(_05639_),
    .Y(_05640_));
 NOR2x1_ASAP7_75t_R _11762_ (.A(net4064),
    .B(net5654),
    .Y(_05641_));
 INVx1_ASAP7_75t_R _11763_ (.A(_05641_),
    .Y(_05642_));
 XOR2x2_ASAP7_75t_R _11764_ (.A(_05640_),
    .B(net3955),
    .Y(_05643_));
 NOR2x1_ASAP7_75t_R _11765_ (.A(net4542),
    .B(_05613_),
    .Y(_05644_));
 AND2x2_ASAP7_75t_R _11766_ (.A(_05613_),
    .B(net4542),
    .Y(_05645_));
 OAI21x1_ASAP7_75t_R _11767_ (.A1(_05644_),
    .A2(_05645_),
    .B(net4456),
    .Y(_05646_));
 INVx1_ASAP7_75t_R _11768_ (.A(net4063),
    .Y(_05647_));
 AOI211x1_ASAP7_75t_R _11769_ (.A1(_05646_),
    .A2(net4344),
    .B(_05647_),
    .C(net3976),
    .Y(_05648_));
 AOI21x1_ASAP7_75t_R _11770_ (.A1(_05637_),
    .A2(_05648_),
    .B(net3992),
    .Y(_05649_));
 AOI21x1_ASAP7_75t_R _11771_ (.A1(_05649_),
    .A2(net3968),
    .B(net3966),
    .Y(_05650_));
 NOR2x1_ASAP7_75t_R _11772_ (.A(net4031),
    .B(net5612),
    .Y(_05651_));
 NOR2x1_ASAP7_75t_R _11773_ (.A(net4065),
    .B(net3938),
    .Y(_05652_));
 OAI21x1_ASAP7_75t_R _11774_ (.A1(_05652_),
    .A2(_05651_),
    .B(net3947),
    .Y(_05653_));
 INVx1_ASAP7_75t_R _11775_ (.A(net4347),
    .Y(_05654_));
 AND3x1_ASAP7_75t_R _11776_ (.A(net4503),
    .B(net4453),
    .C(_05448_),
    .Y(_05655_));
 AND2x2_ASAP7_75t_R _11777_ (.A(_05655_),
    .B(_05568_),
    .Y(_05656_));
 NAND2x1_ASAP7_75t_R _11778_ (.A(_05656_),
    .B(net4394),
    .Y(_05657_));
 OR5x1_ASAP7_75t_R _11779_ (.A(_05657_),
    .B(net4602),
    .C(net4452),
    .D(net4499),
    .E(net4496),
    .Y(_05658_));
 NOR2x1_ASAP7_75t_R _11780_ (.A(_05654_),
    .B(_05658_),
    .Y(_05659_));
 AND2x2_ASAP7_75t_R _11781_ (.A(_05659_),
    .B(net4307),
    .Y(_05660_));
 AO21x1_ASAP7_75t_R _11782_ (.A1(_05660_),
    .A2(net4346),
    .B(net4400),
    .Y(_05661_));
 XOR2x2_ASAP7_75t_R _11783_ (.A(_05661_),
    .B(net4544),
    .Y(_05662_));
 INVx1_ASAP7_75t_R _11784_ (.A(_05662_),
    .Y(_05663_));
 NOR2x1_ASAP7_75t_R _11785_ (.A(net3957),
    .B(net3954),
    .Y(_05664_));
 NOR3x2_ASAP7_75t_R _11786_ (.B(net3992),
    .C(net3938),
    .Y(_05665_),
    .A(_05642_));
 OAI22x1_ASAP7_75t_R _11787_ (.A1(_05653_),
    .A2(net4003),
    .B1(net3946),
    .B2(_05665_),
    .Y(_05666_));
 NOR2x1_ASAP7_75t_R _11788_ (.A(_05643_),
    .B(_05666_),
    .Y(_05667_));
 NOR2x1_ASAP7_75t_R _11789_ (.A(net3992),
    .B(net3939),
    .Y(_05668_));
 OAI21x1_ASAP7_75t_R _11790_ (.A1(net4003),
    .A2(_05653_),
    .B(net3929),
    .Y(_05669_));
 OA21x2_ASAP7_75t_R _11791_ (.A1(_05667_),
    .A2(_05668_),
    .B(_05669_),
    .Y(_05670_));
 NAND2x1_ASAP7_75t_R _11792_ (.A(net4031),
    .B(_05650_),
    .Y(_05671_));
 NAND2x1_ASAP7_75t_R _11793_ (.A(net4065),
    .B(net3938),
    .Y(_05672_));
 AOI21x1_ASAP7_75t_R _11794_ (.A1(_05671_),
    .A2(_05672_),
    .B(net3956),
    .Y(_05673_));
 INVx2_ASAP7_75t_R _11795_ (.A(_05665_),
    .Y(_05674_));
 AOI21x1_ASAP7_75t_R _11796_ (.A1(net4030),
    .A2(_05673_),
    .B(_05674_),
    .Y(_05675_));
 OAI21x1_ASAP7_75t_R _11797_ (.A1(net3946),
    .A2(_05675_),
    .B(net4004),
    .Y(_05676_));
 AOI211x1_ASAP7_75t_R _11798_ (.A1(_05653_),
    .A2(net3929),
    .B(net3946),
    .C(net4003),
    .Y(_05677_));
 INVx1_ASAP7_75t_R _11799_ (.A(_05677_),
    .Y(_05678_));
 NAND2x1_ASAP7_75t_R _11800_ (.A(net3937),
    .B(net3928),
    .Y(_05679_));
 INVx1_ASAP7_75t_R _11801_ (.A(_05679_),
    .Y(_05680_));
 AOI21x1_ASAP7_75t_R _11802_ (.A1(_05676_),
    .A2(_05678_),
    .B(_05680_),
    .Y(_05681_));
 XNOR2x2_ASAP7_75t_R _11803_ (.A(net4397),
    .B(net4189),
    .Y(_05682_));
 INVx1_ASAP7_75t_R _11804_ (.A(_05682_),
    .Y(_05683_));
 INVx1_ASAP7_75t_R _11805_ (.A(_05664_),
    .Y(_05684_));
 NOR2x1_ASAP7_75t_R _11806_ (.A(net4065),
    .B(net4032),
    .Y(_05685_));
 NOR2x1_ASAP7_75t_R _11807_ (.A(_05637_),
    .B(_05638_),
    .Y(_05686_));
 NOR2x1_ASAP7_75t_R _11808_ (.A(_05685_),
    .B(_05686_),
    .Y(_05687_));
 NOR2x1_ASAP7_75t_R _11809_ (.A(_05650_),
    .B(_05687_),
    .Y(_05688_));
 NOR2x1_ASAP7_75t_R _11810_ (.A(net3956),
    .B(net3938),
    .Y(_05689_));
 NOR2x1_ASAP7_75t_R _11811_ (.A(_05689_),
    .B(_05688_),
    .Y(_05690_));
 NAND2x1p5_ASAP7_75t_R _11812_ (.A(_05665_),
    .B(_05690_),
    .Y(_05691_));
 AO21x1_ASAP7_75t_R _11813_ (.A1(_05672_),
    .A2(_05671_),
    .B(_05663_),
    .Y(_05692_));
 AOI21x1_ASAP7_75t_R _11814_ (.A1(_05684_),
    .A2(_05691_),
    .B(_05692_),
    .Y(_05693_));
 INVx1_ASAP7_75t_R _11815_ (.A(net3916),
    .Y(_05694_));
 XOR2x2_ASAP7_75t_R _11816_ (.A(_05693_),
    .B(_05694_),
    .Y(_05695_));
 AO21x1_ASAP7_75t_R _11817_ (.A1(_05681_),
    .A2(net4062),
    .B(_05695_),
    .Y(_05696_));
 AOI22x1_ASAP7_75t_R _11818_ (.A1(_05673_),
    .A2(net4030),
    .B1(_05684_),
    .B2(_05674_),
    .Y(_05697_));
 XOR2x2_ASAP7_75t_R _11819_ (.A(_05697_),
    .B(_05643_),
    .Y(_05698_));
 NAND2x1_ASAP7_75t_R _11820_ (.A(net3895),
    .B(_05696_),
    .Y(_05699_));
 OAI21x1_ASAP7_75t_R _11821_ (.A1(net3884),
    .A2(_05696_),
    .B(_05699_),
    .Y(_05700_));
 INVx1_ASAP7_75t_R _11822_ (.A(_05700_),
    .Y(_05701_));
 NOR2x1p5_ASAP7_75t_R _11823_ (.A(_05698_),
    .B(_05695_),
    .Y(_05702_));
 NAND2x1p5_ASAP7_75t_R _11824_ (.A(_05681_),
    .B(_05683_),
    .Y(_05703_));
 OAI21x1_ASAP7_75t_R _11825_ (.A1(net3884),
    .A2(_05702_),
    .B(_05703_),
    .Y(_05704_));
 XOR2x2_ASAP7_75t_R _11826_ (.A(_05693_),
    .B(net3916),
    .Y(_05705_));
 XOR2x2_ASAP7_75t_R _11827_ (.A(_05704_),
    .B(net3883),
    .Y(_05706_));
 AOI21x1_ASAP7_75t_R _11828_ (.A1(_05702_),
    .A2(_05703_),
    .B(_05670_),
    .Y(_05707_));
 AO21x1_ASAP7_75t_R _11829_ (.A1(_05678_),
    .A2(_05676_),
    .B(net4112),
    .Y(_05708_));
 AO21x1_ASAP7_75t_R _11830_ (.A1(_05669_),
    .A2(_05684_),
    .B(net4004),
    .Y(_05709_));
 AOI21x1_ASAP7_75t_R _11831_ (.A1(net3907),
    .A2(_05709_),
    .B(net3896),
    .Y(_05710_));
 XOR2x2_ASAP7_75t_R _11832_ (.A(_05708_),
    .B(_05710_),
    .Y(_05711_));
 NAND2x1_ASAP7_75t_R _11833_ (.A(_05707_),
    .B(net3880),
    .Y(_05712_));
 OAI21x1_ASAP7_75t_R _11834_ (.A1(_05707_),
    .A2(_05711_),
    .B(_05712_),
    .Y(_05713_));
 NOR2x2_ASAP7_75t_R _11835_ (.A(_05706_),
    .B(_05713_),
    .Y(_05714_));
 AO21x1_ASAP7_75t_R _11836_ (.A1(net4187),
    .A2(net4307),
    .B(net4402),
    .Y(_05715_));
 XOR2x2_ASAP7_75t_R _11837_ (.A(_05715_),
    .B(net4543),
    .Y(_05716_));
 INVx1_ASAP7_75t_R _11838_ (.A(_05670_),
    .Y(_05717_));
 XOR2x2_ASAP7_75t_R _11839_ (.A(_05666_),
    .B(_05643_),
    .Y(_05718_));
 NAND2x1_ASAP7_75t_R _11840_ (.A(_05718_),
    .B(_05705_),
    .Y(_05719_));
 AO21x1_ASAP7_75t_R _11841_ (.A1(_05717_),
    .A2(_05719_),
    .B(net4062),
    .Y(_05720_));
 NAND2x1_ASAP7_75t_R _11842_ (.A(net4062),
    .B(_05707_),
    .Y(_05721_));
 AOI21x1_ASAP7_75t_R _11843_ (.A1(_05684_),
    .A2(_05669_),
    .B(net4030),
    .Y(_05722_));
 NOR2x1_ASAP7_75t_R _11844_ (.A(net3908),
    .B(_05722_),
    .Y(_05723_));
 AOI21x1_ASAP7_75t_R _11845_ (.A1(_05720_),
    .A2(_05721_),
    .B(net3879),
    .Y(_05724_));
 NAND2x1p5_ASAP7_75t_R _11846_ (.A(_05716_),
    .B(_05724_),
    .Y(_05725_));
 OAI21x1_ASAP7_75t_R _11847_ (.A1(_05701_),
    .A2(_05714_),
    .B(_05725_),
    .Y(_05726_));
 XOR2x2_ASAP7_75t_R _11848_ (.A(_05726_),
    .B(net3839),
    .Y(_05727_));
 INVx1_ASAP7_75t_R _11849_ (.A(_05706_),
    .Y(_05728_));
 NOR2x1_ASAP7_75t_R _11850_ (.A(net3839),
    .B(_05726_),
    .Y(_05729_));
 NAND2x1_ASAP7_75t_R _11851_ (.A(net3821),
    .B(net3820),
    .Y(_05730_));
 OAI21x1_ASAP7_75t_R _11852_ (.A1(net3838),
    .A2(_05729_),
    .B(_05730_),
    .Y(_05731_));
 INVx1_ASAP7_75t_R _11853_ (.A(_05731_),
    .Y(_05732_));
 OAI21x1_ASAP7_75t_R _11854_ (.A1(net3908),
    .A2(_05722_),
    .B(net3917),
    .Y(_05733_));
 NOR2x1_ASAP7_75t_R _11855_ (.A(net4112),
    .B(_05733_),
    .Y(_05734_));
 OAI21x1_ASAP7_75t_R _11856_ (.A1(_05719_),
    .A2(_05734_),
    .B(_05717_),
    .Y(_05735_));
 XOR2x2_ASAP7_75t_R _11857_ (.A(_05723_),
    .B(net4112),
    .Y(_05736_));
 NAND2x1_ASAP7_75t_R _11858_ (.A(_05736_),
    .B(_05735_),
    .Y(_05737_));
 OAI21x1_ASAP7_75t_R _11859_ (.A1(net3879),
    .A2(net3863),
    .B(_05737_),
    .Y(_05738_));
 AOI21x1_ASAP7_75t_R _11860_ (.A1(_05714_),
    .A2(_05725_),
    .B(_05701_),
    .Y(_05739_));
 NAND2x1_ASAP7_75t_R _11861_ (.A(net3837),
    .B(_05739_),
    .Y(_05740_));
 INVx1_ASAP7_75t_R _11862_ (.A(_05720_),
    .Y(_05741_));
 NOR2x1_ASAP7_75t_R _11863_ (.A(net4112),
    .B(_05735_),
    .Y(_05742_));
 OAI21x1_ASAP7_75t_R _11864_ (.A1(_05741_),
    .A2(_05742_),
    .B(_05716_),
    .Y(_05743_));
 XNOR2x2_ASAP7_75t_R _11865_ (.A(_05738_),
    .B(_05743_),
    .Y(_05744_));
 NOR2x1_ASAP7_75t_R _11866_ (.A(net3882),
    .B(net5608),
    .Y(_05745_));
 NAND2x1_ASAP7_75t_R _11867_ (.A(net3872),
    .B(_05735_),
    .Y(_05746_));
 OAI21x1_ASAP7_75t_R _11868_ (.A1(net3881),
    .A2(_05745_),
    .B(_05746_),
    .Y(_05747_));
 NAND2x1_ASAP7_75t_R _11869_ (.A(_05728_),
    .B(_05747_),
    .Y(_05748_));
 INVx1_ASAP7_75t_R _11870_ (.A(net4060),
    .Y(_05749_));
 INVx1_ASAP7_75t_R _11871_ (.A(net3879),
    .Y(_05750_));
 OAI21x1_ASAP7_75t_R _11872_ (.A1(_05741_),
    .A2(_05742_),
    .B(_05750_),
    .Y(_05751_));
 NOR2x1_ASAP7_75t_R _11873_ (.A(_05749_),
    .B(_05751_),
    .Y(_05752_));
 OAI21x1_ASAP7_75t_R _11874_ (.A1(_05748_),
    .A2(_05752_),
    .B(net3851),
    .Y(_05753_));
 NAND2x1_ASAP7_75t_R _11875_ (.A(_05744_),
    .B(_05753_),
    .Y(_05754_));
 NAND2x1_ASAP7_75t_R _11876_ (.A(_05754_),
    .B(_05740_),
    .Y(_05755_));
 AO21x1_ASAP7_75t_R _11877_ (.A1(_05748_),
    .A2(net3851),
    .B(net4061),
    .Y(_05756_));
 NAND2x1p5_ASAP7_75t_R _11878_ (.A(_05739_),
    .B(net4061),
    .Y(_05757_));
 AO21x1_ASAP7_75t_R _11879_ (.A1(net4303),
    .A2(net4302),
    .B(net4402),
    .Y(_05758_));
 XNOR2x2_ASAP7_75t_R _11880_ (.A(net4349),
    .B(_05758_),
    .Y(_05759_));
 NAND2x1_ASAP7_75t_R _11881_ (.A(net3864),
    .B(net3850),
    .Y(_05760_));
 INVx1_ASAP7_75t_R _11882_ (.A(_05760_),
    .Y(_05761_));
 NOR2x1_ASAP7_75t_R _11883_ (.A(_05759_),
    .B(_05761_),
    .Y(_05762_));
 INVx1_ASAP7_75t_R _11884_ (.A(_05762_),
    .Y(_05763_));
 AOI21x1_ASAP7_75t_R _11885_ (.A1(_05756_),
    .A2(_05757_),
    .B(_05763_),
    .Y(_05764_));
 NOR2x1p5_ASAP7_75t_R _11886_ (.A(net3781),
    .B(_05755_),
    .Y(_05765_));
 OAI21x1_ASAP7_75t_R _11887_ (.A1(net3798),
    .A2(_05732_),
    .B(_05765_),
    .Y(_05766_));
 OA21x2_ASAP7_75t_R _11888_ (.A1(net3781),
    .A2(net3783),
    .B(_05755_),
    .Y(_05767_));
 INVx1_ASAP7_75t_R _11889_ (.A(_05767_),
    .Y(_05768_));
 NAND2x1_ASAP7_75t_R _11890_ (.A(_05766_),
    .B(_05768_),
    .Y(_05769_));
 INVx1_ASAP7_75t_R _11891_ (.A(net3837),
    .Y(_05770_));
 AOI211x1_ASAP7_75t_R _11892_ (.A1(net3821),
    .A2(net3836),
    .B(net3840),
    .C(_05770_),
    .Y(_05771_));
 XOR2x2_ASAP7_75t_R _11893_ (.A(_05743_),
    .B(_05738_),
    .Y(_05772_));
 NOR2x1_ASAP7_75t_R _11894_ (.A(_05772_),
    .B(net5609),
    .Y(_05773_));
 NOR2x1_ASAP7_75t_R _11895_ (.A(_05771_),
    .B(_05773_),
    .Y(_05774_));
 NAND2x1_ASAP7_75t_R _11896_ (.A(_05727_),
    .B(_05774_),
    .Y(_05775_));
 OAI21x1_ASAP7_75t_R _11897_ (.A1(net5616),
    .A2(_05775_),
    .B(_05731_),
    .Y(_05776_));
 NAND2x1p5_ASAP7_75t_R _11898_ (.A(net3782),
    .B(net5594),
    .Y(_05777_));
 NAND2x1p5_ASAP7_75t_R _11899_ (.A(net3807),
    .B(net3797),
    .Y(_05778_));
 INVx1_ASAP7_75t_R _11900_ (.A(_05778_),
    .Y(_05779_));
 NOR2x1_ASAP7_75t_R _11901_ (.A(net4186),
    .B(_05779_),
    .Y(_05780_));
 INVx1_ASAP7_75t_R _11902_ (.A(_05780_),
    .Y(_05781_));
 INVx1_ASAP7_75t_R _11903_ (.A(_05756_),
    .Y(_05782_));
 AOI211x1_ASAP7_75t_R _11904_ (.A1(net3822),
    .A2(net3834),
    .B(net3841),
    .C(net4029),
    .Y(_05783_));
 OAI21x1_ASAP7_75t_R _11905_ (.A1(_05782_),
    .A2(_05783_),
    .B(net3806),
    .Y(_05784_));
 XOR2x2_ASAP7_75t_R _11906_ (.A(net3809),
    .B(net3835),
    .Y(_05785_));
 NOR2x1_ASAP7_75t_R _11907_ (.A(_05785_),
    .B(_05755_),
    .Y(_05786_));
 AOI21x1_ASAP7_75t_R _11908_ (.A1(_05784_),
    .A2(_05786_),
    .B(_05732_),
    .Y(_05787_));
 NAND2x1_ASAP7_75t_R _11909_ (.A(net4061),
    .B(net3808),
    .Y(_05788_));
 XOR2x2_ASAP7_75t_R _11910_ (.A(_05788_),
    .B(net3819),
    .Y(_05789_));
 INVx1_ASAP7_75t_R _11911_ (.A(_05789_),
    .Y(_05790_));
 OAI21x1_ASAP7_75t_R _11912_ (.A1(_05781_),
    .A2(_05787_),
    .B(_05790_),
    .Y(_05791_));
 NAND2x1_ASAP7_75t_R _11913_ (.A(net3748),
    .B(net3735),
    .Y(_05792_));
 NOR2x1_ASAP7_75t_R _11914_ (.A(net3778),
    .B(_05787_),
    .Y(_05793_));
 AOI21x1_ASAP7_75t_R _11915_ (.A1(_05780_),
    .A2(net5594),
    .B(_05789_),
    .Y(_05794_));
 AOI21x1_ASAP7_75t_R _11916_ (.A1(net3764),
    .A2(net5594),
    .B(net3763),
    .Y(_05795_));
 OAI21x1_ASAP7_75t_R _11917_ (.A1(_05794_),
    .A2(_05793_),
    .B(_05795_),
    .Y(_05796_));
 XOR2x2_ASAP7_75t_R _11918_ (.A(_05766_),
    .B(net3796),
    .Y(_05797_));
 INVx3_ASAP7_75t_R _11919_ (.A(_05797_),
    .Y(_05798_));
 NOR2x1_ASAP7_75t_R _11920_ (.A(net4402),
    .B(net4187),
    .Y(_05799_));
 XNOR2x2_ASAP7_75t_R _11921_ (.A(net4546),
    .B(_05799_),
    .Y(_05800_));
 NAND2x1_ASAP7_75t_R _11922_ (.A(net4186),
    .B(net5593),
    .Y(_05801_));
 INVx1_ASAP7_75t_R _11923_ (.A(net4186),
    .Y(_05802_));
 NAND2x1_ASAP7_75t_R _11924_ (.A(_05787_),
    .B(_05802_),
    .Y(_05803_));
 AOI21x1_ASAP7_75t_R _11925_ (.A1(_05803_),
    .A2(_05801_),
    .B(net3762),
    .Y(_05804_));
 AOI22x1_ASAP7_75t_R _11926_ (.A1(_05796_),
    .A2(_05798_),
    .B1(_05804_),
    .B2(net4059),
    .Y(_05805_));
 NAND2x1_ASAP7_75t_R _11927_ (.A(_05792_),
    .B(_05805_),
    .Y(_05806_));
 AOI21x1_ASAP7_75t_R _11928_ (.A1(net4059),
    .A2(net3733),
    .B(_05796_),
    .Y(_05807_));
 AOI21x1_ASAP7_75t_R _11929_ (.A1(net3749),
    .A2(_05806_),
    .B(_05807_),
    .Y(_05808_));
 INVx1_ASAP7_75t_R _11930_ (.A(_05808_),
    .Y(_05809_));
 INVx1_ASAP7_75t_R _11931_ (.A(_05800_),
    .Y(_05810_));
 NAND3x1_ASAP7_75t_R _11932_ (.A(net3777),
    .B(net3780),
    .C(net3798),
    .Y(_05811_));
 AOI21x1_ASAP7_75t_R _11933_ (.A1(net3783),
    .A2(_05811_),
    .B(_05802_),
    .Y(_05812_));
 NOR2x1p5_ASAP7_75t_R _11934_ (.A(net4186),
    .B(net5593),
    .Y(_05813_));
 OAI21x1_ASAP7_75t_R _11935_ (.A1(_05812_),
    .A2(_05813_),
    .B(net3779),
    .Y(_05814_));
 AOI21x1_ASAP7_75t_R _11936_ (.A1(_05791_),
    .A2(_05777_),
    .B(_05769_),
    .Y(_05815_));
 OAI21x1_ASAP7_75t_R _11937_ (.A1(_05810_),
    .A2(_05814_),
    .B(_05815_),
    .Y(_05816_));
 NAND2x1p5_ASAP7_75t_R _11938_ (.A(net3734),
    .B(_05816_),
    .Y(_05817_));
 OAI21x1_ASAP7_75t_R _11939_ (.A1(_05812_),
    .A2(_05813_),
    .B(_05800_),
    .Y(_05818_));
 NOR2x1_ASAP7_75t_R _11940_ (.A(net3762),
    .B(net5593),
    .Y(_05819_));
 XOR2x2_ASAP7_75t_R _11941_ (.A(_05778_),
    .B(net4186),
    .Y(_05820_));
 NOR2x1_ASAP7_75t_R _11942_ (.A(_05820_),
    .B(_05787_),
    .Y(_05821_));
 NOR2x1_ASAP7_75t_R _11943_ (.A(_05819_),
    .B(_05821_),
    .Y(_05822_));
 XOR2x2_ASAP7_75t_R _11944_ (.A(_05818_),
    .B(_05822_),
    .Y(_05823_));
 AOI211x1_ASAP7_75t_R _11945_ (.A1(_05815_),
    .A2(_05818_),
    .B(net3747),
    .C(net3732),
    .Y(_05824_));
 AOI21x1_ASAP7_75t_R _11946_ (.A1(_05817_),
    .A2(_05823_),
    .B(_05824_),
    .Y(_05825_));
 XOR2x2_ASAP7_75t_R _11947_ (.A(_05805_),
    .B(_05792_),
    .Y(_05826_));
 NAND2x1p5_ASAP7_75t_R _11948_ (.A(_05825_),
    .B(_05826_),
    .Y(_05827_));
 AOI211x1_ASAP7_75t_R _11949_ (.A1(_05815_),
    .A2(_05814_),
    .B(net3747),
    .C(net4028),
    .Y(_05828_));
 AOI21x1_ASAP7_75t_R _11950_ (.A1(net3734),
    .A2(_05816_),
    .B(_05800_),
    .Y(_05829_));
 AO21x1_ASAP7_75t_R _11951_ (.A1(net4391),
    .A2(net4303),
    .B(net4402),
    .Y(_05830_));
 XOR2x2_ASAP7_75t_R _11952_ (.A(_05830_),
    .B(net4398),
    .Y(_05831_));
 INVx1_ASAP7_75t_R _11953_ (.A(_05831_),
    .Y(_05832_));
 NAND2x1_ASAP7_75t_R _11954_ (.A(_05801_),
    .B(_05803_),
    .Y(_05833_));
 INVx1_ASAP7_75t_R _11955_ (.A(_05833_),
    .Y(_05834_));
 NOR2x1_ASAP7_75t_R _11956_ (.A(_05832_),
    .B(_05834_),
    .Y(_05835_));
 OAI21x1_ASAP7_75t_R _11957_ (.A1(_05828_),
    .A2(_05829_),
    .B(_05835_),
    .Y(_05836_));
 INVx2_ASAP7_75t_R _11958_ (.A(_05836_),
    .Y(_05837_));
 AOI21x1_ASAP7_75t_R _11959_ (.A1(_05809_),
    .A2(net5939),
    .B(_05837_),
    .Y(_05838_));
 XOR2x2_ASAP7_75t_R _11960_ (.A(_05838_),
    .B(net3681),
    .Y(_05839_));
 XOR2x2_ASAP7_75t_R _11961_ (.A(_05833_),
    .B(net4027),
    .Y(_05840_));
 AO21x1_ASAP7_75t_R _11962_ (.A1(_05816_),
    .A2(net3734),
    .B(_05840_),
    .Y(_05841_));
 OAI21x1_ASAP7_75t_R _11963_ (.A1(net3716),
    .A2(net3694),
    .B(_05841_),
    .Y(_05842_));
 INVx1_ASAP7_75t_R _11964_ (.A(net3679),
    .Y(_05843_));
 OAI21x1_ASAP7_75t_R _11965_ (.A1(_05827_),
    .A2(_05837_),
    .B(_05809_),
    .Y(_05844_));
 NOR2x1_ASAP7_75t_R _11966_ (.A(_05844_),
    .B(_05843_),
    .Y(_05845_));
 OAI21x1_ASAP7_75t_R _11967_ (.A1(net3707),
    .A2(net3693),
    .B(net4185),
    .Y(_05846_));
 XOR2x2_ASAP7_75t_R _11968_ (.A(_05842_),
    .B(_05846_),
    .Y(_05847_));
 INVx1_ASAP7_75t_R _11969_ (.A(_05824_),
    .Y(_05848_));
 OAI21x1_ASAP7_75t_R _11970_ (.A1(net3747),
    .A2(_05807_),
    .B(_05823_),
    .Y(_05849_));
 NAND2x1_ASAP7_75t_R _11971_ (.A(_05848_),
    .B(_05849_),
    .Y(_05850_));
 XNOR2x2_ASAP7_75t_R _11972_ (.A(_05792_),
    .B(_05805_),
    .Y(_05851_));
 NOR2x1_ASAP7_75t_R _11973_ (.A(_05850_),
    .B(_05851_),
    .Y(_05852_));
 AOI21x1_ASAP7_75t_R _11974_ (.A1(net5599),
    .A2(_05852_),
    .B(net3695),
    .Y(_05853_));
 NOR2x1_ASAP7_75t_R _11975_ (.A(_05847_),
    .B(_05853_),
    .Y(_05854_));
 NOR2x1_ASAP7_75t_R _11976_ (.A(_05854_),
    .B(_05845_),
    .Y(_05855_));
 NAND2x1_ASAP7_75t_R _11977_ (.A(_05855_),
    .B(_05839_),
    .Y(_05856_));
 INVx1_ASAP7_75t_R _11978_ (.A(net3707),
    .Y(_05857_));
 INVx1_ASAP7_75t_R _11979_ (.A(net3693),
    .Y(_05858_));
 NAND2x1_ASAP7_75t_R _11980_ (.A(_05857_),
    .B(_05858_),
    .Y(_05859_));
 INVx1_ASAP7_75t_R _11981_ (.A(_05859_),
    .Y(_05860_));
 NAND3x1_ASAP7_75t_R _11982_ (.A(net3680),
    .B(net3708),
    .C(net3681),
    .Y(_05861_));
 AOI21x1_ASAP7_75t_R _11983_ (.A1(net3682),
    .A2(_05861_),
    .B(net4185),
    .Y(_05862_));
 NOR2x1_ASAP7_75t_R _11984_ (.A(net4111),
    .B(_05844_),
    .Y(_05863_));
 NAND2x1_ASAP7_75t_R _11985_ (.A(net4456),
    .B(net4249),
    .Y(_05864_));
 XOR2x2_ASAP7_75t_R _11986_ (.A(_05864_),
    .B(net4601),
    .Y(_05865_));
 OAI21x1_ASAP7_75t_R _11987_ (.A1(_05863_),
    .A2(_05862_),
    .B(net4109),
    .Y(_05866_));
 NOR2x1p5_ASAP7_75t_R _11988_ (.A(_05860_),
    .B(_05866_),
    .Y(_05867_));
 NOR2x1_ASAP7_75t_R _11989_ (.A(net3602),
    .B(net3601),
    .Y(_05868_));
 NAND2x1p5_ASAP7_75t_R _11990_ (.A(net4111),
    .B(_05844_),
    .Y(_05869_));
 NAND2x1_ASAP7_75t_R _11991_ (.A(net4185),
    .B(_05853_),
    .Y(_05870_));
 INVx1_ASAP7_75t_R _11992_ (.A(_05865_),
    .Y(_05871_));
 AOI21x1_ASAP7_75t_R _11993_ (.A1(_05869_),
    .A2(_05870_),
    .B(_05871_),
    .Y(_05872_));
 NAND2x1_ASAP7_75t_R _11994_ (.A(net3679),
    .B(_05853_),
    .Y(_05873_));
 OAI21x1_ASAP7_75t_R _11995_ (.A1(_05853_),
    .A2(net3665),
    .B(_05873_),
    .Y(_05874_));
 AO21x1_ASAP7_75t_R _11996_ (.A1(_05872_),
    .A2(net3664),
    .B(_05874_),
    .Y(_05875_));
 NAND2x1_ASAP7_75t_R _11997_ (.A(net3681),
    .B(_05838_),
    .Y(_05876_));
 INVx1_ASAP7_75t_R _11998_ (.A(_05861_),
    .Y(_05877_));
 AO21x1_ASAP7_75t_R _11999_ (.A1(_05876_),
    .A2(net3706),
    .B(_05877_),
    .Y(_05878_));
 XOR2x2_ASAP7_75t_R _12000_ (.A(net3678),
    .B(_05838_),
    .Y(_05879_));
 OA21x2_ASAP7_75t_R _12001_ (.A1(_05875_),
    .A2(net3622),
    .B(_05879_),
    .Y(_05880_));
 NOR2x1p5_ASAP7_75t_R _12002_ (.A(_05868_),
    .B(_05880_),
    .Y(_05881_));
 INVx1_ASAP7_75t_R _12003_ (.A(_05878_),
    .Y(_05882_));
 NOR2x1_ASAP7_75t_R _12004_ (.A(_05879_),
    .B(_05874_),
    .Y(_05883_));
 NAND2x1_ASAP7_75t_R _12005_ (.A(net3664),
    .B(_05872_),
    .Y(_05884_));
 OAI21x1_ASAP7_75t_R _12006_ (.A1(_05882_),
    .A2(_05883_),
    .B(_05884_),
    .Y(_05885_));
 XOR2x2_ASAP7_75t_R _12007_ (.A(_05885_),
    .B(net3624),
    .Y(_05886_));
 NOR2x1_ASAP7_75t_R _12008_ (.A(_05886_),
    .B(_05881_),
    .Y(_05887_));
 NOR2x1_ASAP7_75t_R _12009_ (.A(net4303),
    .B(net4402),
    .Y(_05888_));
 XOR2x2_ASAP7_75t_R _12010_ (.A(_05888_),
    .B(net4399),
    .Y(_05889_));
 OAI21x1_ASAP7_75t_R _12011_ (.A1(_05867_),
    .A2(_05856_),
    .B(net3622),
    .Y(_05890_));
 NAND2x1p5_ASAP7_75t_R _12012_ (.A(_05890_),
    .B(net4058),
    .Y(_05891_));
 AOI21x1_ASAP7_75t_R _12013_ (.A1(_05884_),
    .A2(_05883_),
    .B(_05882_),
    .Y(_05892_));
 NAND2x1_ASAP7_75t_R _12014_ (.A(_05892_),
    .B(net4110),
    .Y(_05893_));
 NAND2x1_ASAP7_75t_R _12015_ (.A(net3644),
    .B(net3643),
    .Y(_05894_));
 INVx1_ASAP7_75t_R _12016_ (.A(_05894_),
    .Y(_05895_));
 AOI21x1_ASAP7_75t_R _12017_ (.A1(_05891_),
    .A2(_05893_),
    .B(_05895_),
    .Y(_05896_));
 XOR2x2_ASAP7_75t_R _12018_ (.A(_05859_),
    .B(net4185),
    .Y(_05897_));
 NOR2x1_ASAP7_75t_R _12019_ (.A(_05860_),
    .B(_05844_),
    .Y(_05898_));
 AO21x1_ASAP7_75t_R _12020_ (.A1(_05844_),
    .A2(_05897_),
    .B(_05898_),
    .Y(_05899_));
 XOR2x2_ASAP7_75t_R _12021_ (.A(_05899_),
    .B(net3623),
    .Y(_05900_));
 NAND2x1_ASAP7_75t_R _12022_ (.A(net3620),
    .B(_05892_),
    .Y(_05901_));
 OAI21x1_ASAP7_75t_R _12023_ (.A1(_05892_),
    .A2(_05900_),
    .B(_05901_),
    .Y(_05902_));
 AOI21x1_ASAP7_75t_R _12024_ (.A1(_05896_),
    .A2(net4184),
    .B(_05902_),
    .Y(_05903_));
 OAI21x1_ASAP7_75t_R _12025_ (.A1(net3588),
    .A2(_05887_),
    .B(_05903_),
    .Y(_05904_));
 XOR2x2_ASAP7_75t_R _12026_ (.A(net3587),
    .B(_05904_),
    .Y(_05905_));
 INVx3_ASAP7_75t_R _12027_ (.A(_05905_),
    .Y(_05906_));
 INVx1_ASAP7_75t_R _12028_ (.A(_05881_),
    .Y(_05907_));
 INVx1_ASAP7_75t_R _12029_ (.A(_05889_),
    .Y(_05908_));
 NOR2x1_ASAP7_75t_R _12030_ (.A(net4058),
    .B(_05890_),
    .Y(_05909_));
 NOR2x1_ASAP7_75t_R _12031_ (.A(net4110),
    .B(_05892_),
    .Y(_05910_));
 OAI21x1_ASAP7_75t_R _12032_ (.A1(_05909_),
    .A2(_05910_),
    .B(net3621),
    .Y(_05911_));
 NOR2x1p5_ASAP7_75t_R _12033_ (.A(net4108),
    .B(_05911_),
    .Y(_05912_));
 OAI21x1_ASAP7_75t_R _12034_ (.A1(_05907_),
    .A2(net3556),
    .B(net3570),
    .Y(_05913_));
 NAND2x1_ASAP7_75t_R _12035_ (.A(_05913_),
    .B(_05904_),
    .Y(_05914_));
 NAND2x1_ASAP7_75t_R _12036_ (.A(_05657_),
    .B(net4456),
    .Y(_05915_));
 OA21x2_ASAP7_75t_R _12037_ (.A1(net4400),
    .A2(net4451),
    .B(_05915_),
    .Y(_05916_));
 XOR2x2_ASAP7_75t_R _12038_ (.A(_05916_),
    .B(net4496),
    .Y(_05917_));
 INVx1_ASAP7_75t_R _12039_ (.A(_05917_),
    .Y(_05918_));
 NOR2x1_ASAP7_75t_R _12040_ (.A(_05902_),
    .B(_05886_),
    .Y(_05919_));
 NAND2x1_ASAP7_75t_R _12041_ (.A(net4184),
    .B(_05896_),
    .Y(_05920_));
 AOI21x1_ASAP7_75t_R _12042_ (.A1(_05919_),
    .A2(_05920_),
    .B(net3588),
    .Y(_05921_));
 NOR2x1_ASAP7_75t_R _12043_ (.A(net4184),
    .B(_05921_),
    .Y(_05922_));
 NAND2x1_ASAP7_75t_R _12044_ (.A(_05900_),
    .B(_05890_),
    .Y(_05923_));
 OAI21x1_ASAP7_75t_R _12045_ (.A1(net3620),
    .A2(net5595),
    .B(_05923_),
    .Y(_05924_));
 INVx1_ASAP7_75t_R _12046_ (.A(_05886_),
    .Y(_05925_));
 NAND2x1_ASAP7_75t_R _12047_ (.A(_05924_),
    .B(_05925_),
    .Y(_05926_));
 OAI21x1_ASAP7_75t_R _12048_ (.A1(_05926_),
    .A2(_05912_),
    .B(_05907_),
    .Y(_05927_));
 NOR2x1_ASAP7_75t_R _12049_ (.A(net4108),
    .B(_05927_),
    .Y(_05928_));
 NAND2x1_ASAP7_75t_R _12050_ (.A(net3586),
    .B(net3585),
    .Y(_05929_));
 OAI21x1_ASAP7_75t_R _12051_ (.A1(_05928_),
    .A2(_05922_),
    .B(_05929_),
    .Y(_05930_));
 AO21x2_ASAP7_75t_R _12052_ (.A1(_05893_),
    .A2(_05891_),
    .B(_05908_),
    .Y(_05931_));
 INVx1_ASAP7_75t_R _12053_ (.A(_05931_),
    .Y(_05932_));
 NAND2x1_ASAP7_75t_R _12054_ (.A(_05890_),
    .B(net4110),
    .Y(_05933_));
 XOR2x2_ASAP7_75t_R _12055_ (.A(_05933_),
    .B(_05895_),
    .Y(_05934_));
 AND3x4_ASAP7_75t_R _12056_ (.A(_05932_),
    .B(_05934_),
    .C(net3588),
    .Y(_05935_));
 OAI21x1_ASAP7_75t_R _12057_ (.A1(_05934_),
    .A2(_05926_),
    .B(_05907_),
    .Y(_05936_));
 AOI21x1_ASAP7_75t_R _12058_ (.A1(net3554),
    .A2(_05936_),
    .B(net3567),
    .Y(_05937_));
 NOR2x1_ASAP7_75t_R _12059_ (.A(_05935_),
    .B(_05937_),
    .Y(_05938_));
 INVx1_ASAP7_75t_R _12060_ (.A(_05938_),
    .Y(_05939_));
 OAI21x1_ASAP7_75t_R _12061_ (.A1(_05918_),
    .A2(_05930_),
    .B(_05939_),
    .Y(_05940_));
 AOI21x1_ASAP7_75t_R _12062_ (.A1(_05906_),
    .A2(net3527),
    .B(_05940_),
    .Y(_05941_));
 AOI21x1_ASAP7_75t_R _12063_ (.A1(net3588),
    .A2(net3555),
    .B(net3569),
    .Y(_05942_));
 AOI21x1_ASAP7_75t_R _12064_ (.A1(net3557),
    .A2(net3544),
    .B(_05942_),
    .Y(_05943_));
 XOR2x2_ASAP7_75t_R _12065_ (.A(_05941_),
    .B(net3525),
    .Y(_05944_));
 NAND2x1_ASAP7_75t_R _12066_ (.A(net4108),
    .B(net3544),
    .Y(_05945_));
 NAND2x1_ASAP7_75t_R _12067_ (.A(net4184),
    .B(net3545),
    .Y(_05946_));
 AO21x1_ASAP7_75t_R _12068_ (.A1(_05945_),
    .A2(_05946_),
    .B(_05918_),
    .Y(_05947_));
 INVx2_ASAP7_75t_R _12069_ (.A(_05935_),
    .Y(_05948_));
 XOR2x2_ASAP7_75t_R _12070_ (.A(net5610),
    .B(net3621),
    .Y(_05949_));
 AOI21x1_ASAP7_75t_R _12071_ (.A1(_05949_),
    .A2(_05919_),
    .B(net3588),
    .Y(_05950_));
 OAI21x1_ASAP7_75t_R _12072_ (.A1(_05931_),
    .A2(_05950_),
    .B(_05949_),
    .Y(_05951_));
 AOI21x1_ASAP7_75t_R _12073_ (.A1(_05951_),
    .A2(_05948_),
    .B(_05914_),
    .Y(_05952_));
 INVx1_ASAP7_75t_R _12074_ (.A(net3568),
    .Y(_05953_));
 AOI21x1_ASAP7_75t_R _12075_ (.A1(_05946_),
    .A2(_05945_),
    .B(_05953_),
    .Y(_05954_));
 NAND2x1_ASAP7_75t_R _12076_ (.A(net4107),
    .B(_05954_),
    .Y(_05955_));
 AOI21x1_ASAP7_75t_R _12077_ (.A1(net3508),
    .A2(_05955_),
    .B(net3528),
    .Y(_05956_));
 NAND2x1_ASAP7_75t_R _12078_ (.A(net3554),
    .B(net3542),
    .Y(_05957_));
 AO21x1_ASAP7_75t_R _12079_ (.A1(net3544),
    .A2(net4184),
    .B(net3568),
    .Y(_05958_));
 NAND2x1_ASAP7_75t_R _12080_ (.A(_05957_),
    .B(_05958_),
    .Y(_05959_));
 OAI21x1_ASAP7_75t_R _12081_ (.A1(net3509),
    .A2(_05956_),
    .B(net3507),
    .Y(_05960_));
 INVx1_ASAP7_75t_R _12082_ (.A(_05959_),
    .Y(_05961_));
 OAI21x1_ASAP7_75t_R _12083_ (.A1(_05930_),
    .A2(_05918_),
    .B(_05952_),
    .Y(_05962_));
 AOI21x1_ASAP7_75t_R _12084_ (.A1(_05906_),
    .A2(_05962_),
    .B(_05947_),
    .Y(_05963_));
 NAND2x1_ASAP7_75t_R _12085_ (.A(_05961_),
    .B(_05963_),
    .Y(_05964_));
 NOR2x1_ASAP7_75t_R _12086_ (.A(_05918_),
    .B(_05930_),
    .Y(_05965_));
 OAI21x1_ASAP7_75t_R _12087_ (.A1(_05965_),
    .A2(_05906_),
    .B(net3510),
    .Y(_05966_));
 OAI21x1_ASAP7_75t_R _12088_ (.A1(net3488),
    .A2(_05956_),
    .B(net5941),
    .Y(_05967_));
 AOI21x1_ASAP7_75t_R _12089_ (.A1(_05960_),
    .A2(_05964_),
    .B(_05967_),
    .Y(_05968_));
 NAND2x1_ASAP7_75t_R _12090_ (.A(net3523),
    .B(net3524),
    .Y(_05969_));
 OAI21x1_ASAP7_75t_R _12091_ (.A1(net3543),
    .A2(net3526),
    .B(_05943_),
    .Y(_05970_));
 NOR2x1_ASAP7_75t_R _12092_ (.A(_05930_),
    .B(_05970_),
    .Y(_05971_));
 OAI21x1_ASAP7_75t_R _12093_ (.A1(_05954_),
    .A2(_05970_),
    .B(net3511),
    .Y(_05972_));
 OAI21x1_ASAP7_75t_R _12094_ (.A1(_05971_),
    .A2(_05972_),
    .B(net4057),
    .Y(_05973_));
 AOI211x1_ASAP7_75t_R _12095_ (.A1(_05930_),
    .A2(_05952_),
    .B(net3528),
    .C(_05918_),
    .Y(_05974_));
 INVx1_ASAP7_75t_R _12096_ (.A(_05974_),
    .Y(_05975_));
 AOI211x1_ASAP7_75t_R _12097_ (.A1(net4345),
    .A2(_05584_),
    .B(net4504),
    .C(net4506),
    .Y(_05976_));
 XNOR2x2_ASAP7_75t_R _12098_ (.A(net4499),
    .B(_05976_),
    .Y(_05977_));
 INVx1_ASAP7_75t_R _12099_ (.A(_05977_),
    .Y(_05978_));
 AOI21x1_ASAP7_75t_R _12100_ (.A1(_05973_),
    .A2(_05975_),
    .B(_05978_),
    .Y(_05979_));
 NAND2x1_ASAP7_75t_R _12101_ (.A(_05969_),
    .B(_05979_),
    .Y(_05980_));
 OAI21x1_ASAP7_75t_R _12102_ (.A1(net3468),
    .A2(_05968_),
    .B(_05980_),
    .Y(_05981_));
 NAND2x1_ASAP7_75t_R _12103_ (.A(net3479),
    .B(net3478),
    .Y(_05982_));
 XOR2x2_ASAP7_75t_R _12104_ (.A(_05981_),
    .B(_05982_),
    .Y(_05983_));
 AOI21x1_ASAP7_75t_R _12105_ (.A1(net3512),
    .A2(_05962_),
    .B(net4057),
    .Y(_05984_));
 INVx1_ASAP7_75t_R _12106_ (.A(_05963_),
    .Y(_05985_));
 OAI21x1_ASAP7_75t_R _12107_ (.A1(_05969_),
    .A2(_05984_),
    .B(_05985_),
    .Y(_05986_));
 AOI21x1_ASAP7_75t_R _12108_ (.A1(net3512),
    .A2(_05962_),
    .B(net4107),
    .Y(_05987_));
 OAI21x1_ASAP7_75t_R _12109_ (.A1(_05974_),
    .A2(_05987_),
    .B(_05977_),
    .Y(_05988_));
 XOR2x2_ASAP7_75t_R _12110_ (.A(_05986_),
    .B(_05988_),
    .Y(_05989_));
 INVx1_ASAP7_75t_R _12111_ (.A(_05969_),
    .Y(_05990_));
 NOR2x1_ASAP7_75t_R _12112_ (.A(_05990_),
    .B(_05988_),
    .Y(_05991_));
 NOR2x1_ASAP7_75t_R _12113_ (.A(_05963_),
    .B(_05961_),
    .Y(_05992_));
 AOI211x1_ASAP7_75t_R _12114_ (.A1(net3493),
    .A2(net3513),
    .B(net3509),
    .C(net3507),
    .Y(_05993_));
 INVx1_ASAP7_75t_R _12115_ (.A(_05966_),
    .Y(_05994_));
 NOR2x1_ASAP7_75t_R _12116_ (.A(_05994_),
    .B(_05941_),
    .Y(_05995_));
 OAI21x1_ASAP7_75t_R _12117_ (.A1(_05992_),
    .A2(_05993_),
    .B(_05995_),
    .Y(_05996_));
 INVx1_ASAP7_75t_R _12118_ (.A(_05944_),
    .Y(_05997_));
 OAI21x1_ASAP7_75t_R _12119_ (.A1(_05996_),
    .A2(_05991_),
    .B(_05997_),
    .Y(_05998_));
 NAND2x1_ASAP7_75t_R _12120_ (.A(_05989_),
    .B(_05998_),
    .Y(_05999_));
 INVx1_ASAP7_75t_R _12121_ (.A(_05986_),
    .Y(_06000_));
 AOI21x1_ASAP7_75t_R _12122_ (.A1(_05968_),
    .A2(_05980_),
    .B(_05944_),
    .Y(_06001_));
 NAND2x1_ASAP7_75t_R _12123_ (.A(_06000_),
    .B(_06001_),
    .Y(_06002_));
 NAND2x1p5_ASAP7_75t_R _12124_ (.A(_05999_),
    .B(_06002_),
    .Y(_06003_));
 NOR2x2_ASAP7_75t_R _12125_ (.A(_05983_),
    .B(_06003_),
    .Y(_06004_));
 INVx1_ASAP7_75t_R _12126_ (.A(_06004_),
    .Y(_06005_));
 XOR2x2_ASAP7_75t_R _12127_ (.A(net4248),
    .B(net4602),
    .Y(_06006_));
 INVx1_ASAP7_75t_R _12128_ (.A(_06006_),
    .Y(_06007_));
 NOR2x1_ASAP7_75t_R _12129_ (.A(net4183),
    .B(_05998_),
    .Y(_06008_));
 NOR2x1_ASAP7_75t_R _12130_ (.A(net4247),
    .B(net3451),
    .Y(_06009_));
 NAND2x1_ASAP7_75t_R _12131_ (.A(net3487),
    .B(net3486),
    .Y(_06010_));
 OAI21x1_ASAP7_75t_R _12132_ (.A1(_06008_),
    .A2(_06009_),
    .B(net3477),
    .Y(_06011_));
 NOR2x1_ASAP7_75t_R _12133_ (.A(_06007_),
    .B(_06011_),
    .Y(_06012_));
 INVx1_ASAP7_75t_R _12134_ (.A(_05982_),
    .Y(_06013_));
 NOR2x1_ASAP7_75t_R _12135_ (.A(_06013_),
    .B(net3453),
    .Y(_06014_));
 NOR2x1_ASAP7_75t_R _12136_ (.A(net3467),
    .B(net3452),
    .Y(_06015_));
 INVx1_ASAP7_75t_R _12137_ (.A(_06015_),
    .Y(_06016_));
 OA21x2_ASAP7_75t_R _12138_ (.A1(_06014_),
    .A2(net3466),
    .B(_06016_),
    .Y(_06017_));
 BUFx3_ASAP7_75t_R place2939 (.A(_06311_),
    .Y(net2939));
 INVx1_ASAP7_75t_R _12140_ (.A(_06017_),
    .Y(_06019_));
 OAI21x1_ASAP7_75t_R _12141_ (.A1(_06005_),
    .A2(_06012_),
    .B(_06019_),
    .Y(_06020_));
 NAND2x1p5_ASAP7_75t_R _12142_ (.A(_05998_),
    .B(net4183),
    .Y(_06021_));
 NAND2x1_ASAP7_75t_R _12143_ (.A(net4247),
    .B(_06001_),
    .Y(_06022_));
 INVx1_ASAP7_75t_R _12144_ (.A(_06010_),
    .Y(_06023_));
 AOI21x1_ASAP7_75t_R _12145_ (.A1(_06021_),
    .A2(_06022_),
    .B(_06023_),
    .Y(_06024_));
 NAND2x2_ASAP7_75t_R _12146_ (.A(_06024_),
    .B(_06006_),
    .Y(_06025_));
 XOR2x2_ASAP7_75t_R _12147_ (.A(_06025_),
    .B(net3409),
    .Y(_06026_));
 INVx1_ASAP7_75t_R _12148_ (.A(net3409),
    .Y(_06027_));
 NOR2x1_ASAP7_75t_R _12149_ (.A(_06027_),
    .B(_06017_),
    .Y(_06028_));
 AOI21x1_ASAP7_75t_R _12150_ (.A1(_06020_),
    .A2(_06026_),
    .B(_06028_),
    .Y(_06029_));
 INVx1_ASAP7_75t_R _12151_ (.A(_06029_),
    .Y(_06030_));
 OAI21x1_ASAP7_75t_R _12152_ (.A1(_06008_),
    .A2(_06009_),
    .B(_06006_),
    .Y(_06031_));
 XOR2x2_ASAP7_75t_R _12153_ (.A(_06010_),
    .B(net4247),
    .Y(_06032_));
 NAND2x1_ASAP7_75t_R _12154_ (.A(_06032_),
    .B(net3433),
    .Y(_06033_));
 OAI21x1_ASAP7_75t_R _12155_ (.A1(net3465),
    .A2(net3433),
    .B(_06033_),
    .Y(_06034_));
 INVx1_ASAP7_75t_R _12156_ (.A(_06034_),
    .Y(_06035_));
 AOI211x1_ASAP7_75t_R _12157_ (.A1(_06004_),
    .A2(_06031_),
    .B(_06035_),
    .C(net3408),
    .Y(_06036_));
 XOR2x2_ASAP7_75t_R _12158_ (.A(_06031_),
    .B(_06034_),
    .Y(_06037_));
 AOI21x1_ASAP7_75t_R _12159_ (.A1(_06025_),
    .A2(_06004_),
    .B(_06017_),
    .Y(_06038_));
 NOR2x1_ASAP7_75t_R _12160_ (.A(_06038_),
    .B(_06037_),
    .Y(_06039_));
 NOR2x1p5_ASAP7_75t_R _12161_ (.A(net5632),
    .B(_06039_),
    .Y(_06040_));
 NAND2x2_ASAP7_75t_R _12162_ (.A(_06004_),
    .B(_06025_),
    .Y(_06041_));
 OAI21x1_ASAP7_75t_R _12163_ (.A1(_06007_),
    .A2(_06011_),
    .B(_06027_),
    .Y(_06042_));
 OAI21x1_ASAP7_75t_R _12164_ (.A1(_06019_),
    .A2(_06042_),
    .B(net3434),
    .Y(_06043_));
 NAND2x1_ASAP7_75t_R _12165_ (.A(_06041_),
    .B(_06043_),
    .Y(_06044_));
 NAND2x1p5_ASAP7_75t_R _12166_ (.A(_06040_),
    .B(net5628),
    .Y(_06045_));
 NOR2x1_ASAP7_75t_R _12167_ (.A(net4345),
    .B(net4400),
    .Y(_06046_));
 INVx1_ASAP7_75t_R _12168_ (.A(_05557_),
    .Y(_06047_));
 XOR2x2_ASAP7_75t_R _12169_ (.A(_06046_),
    .B(_06047_),
    .Y(_06048_));
 INVx1_ASAP7_75t_R _12170_ (.A(net4245),
    .Y(_06049_));
 OA21x2_ASAP7_75t_R _12171_ (.A1(_06004_),
    .A2(_06017_),
    .B(net4106),
    .Y(_06050_));
 AOI211x1_ASAP7_75t_R _12172_ (.A1(_06004_),
    .A2(_06011_),
    .B(_06017_),
    .C(net4106),
    .Y(_06051_));
 NAND2x1_ASAP7_75t_R _12173_ (.A(net3419),
    .B(net3431),
    .Y(_06052_));
 OAI21x1_ASAP7_75t_R _12174_ (.A1(_06050_),
    .A2(net5601),
    .B(net3406),
    .Y(_06053_));
 NOR2x1_ASAP7_75t_R _12175_ (.A(_06053_),
    .B(_06049_),
    .Y(_06054_));
 AOI21x1_ASAP7_75t_R _12176_ (.A1(net3358),
    .A2(_06045_),
    .B(net5624),
    .Y(_06055_));
 NAND2x1_ASAP7_75t_R _12177_ (.A(net3359),
    .B(_06055_),
    .Y(_06056_));
 NOR2x1_ASAP7_75t_R _12178_ (.A(net3340),
    .B(net3357),
    .Y(_06057_));
 AOI21x1_ASAP7_75t_R _12179_ (.A1(net3341),
    .A2(_06056_),
    .B(_06057_),
    .Y(_06058_));
 NAND2x1_ASAP7_75t_R _12180_ (.A(net3406),
    .B(_06038_),
    .Y(_06059_));
 XOR2x2_ASAP7_75t_R _12181_ (.A(_06052_),
    .B(_06007_),
    .Y(_06060_));
 NOR2x1p5_ASAP7_75t_R _12182_ (.A(_06060_),
    .B(_06038_),
    .Y(_06061_));
 INVx2_ASAP7_75t_R _12183_ (.A(_06061_),
    .Y(_06062_));
 NAND2x1p5_ASAP7_75t_R _12184_ (.A(net5631),
    .B(_06062_),
    .Y(_06063_));
 OAI21x1_ASAP7_75t_R _12185_ (.A1(_06050_),
    .A2(_06051_),
    .B(_06048_),
    .Y(_06064_));
 XOR2x2_ASAP7_75t_R _12186_ (.A(_06063_),
    .B(net3369),
    .Y(_06065_));
 INVx1_ASAP7_75t_R _12187_ (.A(_06036_),
    .Y(_06066_));
 OAI21x1_ASAP7_75t_R _12188_ (.A1(net5596),
    .A2(net3393),
    .B(_06066_),
    .Y(_06067_));
 OAI21x1_ASAP7_75t_R _12189_ (.A1(_06067_),
    .A2(_06030_),
    .B(_06044_),
    .Y(_06068_));
 INVx1_ASAP7_75t_R _12190_ (.A(_06064_),
    .Y(_06069_));
 INVx1_ASAP7_75t_R _12191_ (.A(_06041_),
    .Y(_06070_));
 AOI21x1_ASAP7_75t_R _12192_ (.A1(net4182),
    .A2(net3407),
    .B(net3409),
    .Y(_06071_));
 INVx1_ASAP7_75t_R _12193_ (.A(net3434),
    .Y(_06072_));
 AOI21x1_ASAP7_75t_R _12194_ (.A1(net3408),
    .A2(_06071_),
    .B(_06072_),
    .Y(_06073_));
 NOR2x1_ASAP7_75t_R _12195_ (.A(_06070_),
    .B(_06073_),
    .Y(_06074_));
 AOI21x1_ASAP7_75t_R _12196_ (.A1(_06059_),
    .A2(_06062_),
    .B(_06074_),
    .Y(_06075_));
 NAND2x1_ASAP7_75t_R _12197_ (.A(_06075_),
    .B(_06069_),
    .Y(_06076_));
 NAND2x1p5_ASAP7_75t_R _12198_ (.A(_06068_),
    .B(_06076_),
    .Y(_06077_));
 AOI21x1_ASAP7_75t_R _12199_ (.A1(net5628),
    .A2(_06040_),
    .B(_06074_),
    .Y(_06078_));
 NOR2x1_ASAP7_75t_R _12200_ (.A(net3420),
    .B(net3432),
    .Y(_06079_));
 NOR2x1_ASAP7_75t_R _12201_ (.A(_06079_),
    .B(_06020_),
    .Y(_06080_));
 OAI21x1_ASAP7_75t_R _12202_ (.A1(net5630),
    .A2(_06080_),
    .B(_06044_),
    .Y(_06081_));
 NOR2x1_ASAP7_75t_R _12203_ (.A(_06064_),
    .B(_06081_),
    .Y(_06082_));
 OAI21x1_ASAP7_75t_R _12204_ (.A1(_06078_),
    .A2(_06082_),
    .B(net3339),
    .Y(_06083_));
 OAI21x1_ASAP7_75t_R _12205_ (.A1(_06065_),
    .A2(_06077_),
    .B(_06083_),
    .Y(_06084_));
 XOR2x2_ASAP7_75t_R _12206_ (.A(_06067_),
    .B(_06054_),
    .Y(_06085_));
 OAI21x1_ASAP7_75t_R _12207_ (.A1(_06078_),
    .A2(_06082_),
    .B(net3356),
    .Y(_06086_));
 OAI21x1_ASAP7_75t_R _12208_ (.A1(_06077_),
    .A2(_06085_),
    .B(_06086_),
    .Y(_06087_));
 NOR2x1p5_ASAP7_75t_R _12209_ (.A(_06084_),
    .B(_06087_),
    .Y(_06088_));
 NOR2x1_ASAP7_75t_R _12210_ (.A(net3380),
    .B(net3379),
    .Y(_06089_));
 INVx1_ASAP7_75t_R _12211_ (.A(_06089_),
    .Y(_06090_));
 AO21x2_ASAP7_75t_R _12212_ (.A1(_06045_),
    .A2(net3358),
    .B(net4246),
    .Y(_06091_));
 OAI21x1_ASAP7_75t_R _12213_ (.A1(_06078_),
    .A2(_06082_),
    .B(net4246),
    .Y(_06092_));
 NOR2x1_ASAP7_75t_R _12214_ (.A(net4343),
    .B(net4400),
    .Y(_06093_));
 XOR2x2_ASAP7_75t_R _12215_ (.A(_06093_),
    .B(net4392),
    .Y(_06094_));
 INVx1_ASAP7_75t_R _12216_ (.A(_06094_),
    .Y(_06095_));
 AOI21x1_ASAP7_75t_R _12217_ (.A1(_06091_),
    .A2(_06092_),
    .B(_06095_),
    .Y(_06096_));
 NAND2x1p5_ASAP7_75t_R _12218_ (.A(_06096_),
    .B(_06090_),
    .Y(_06097_));
 OAI21x1_ASAP7_75t_R _12219_ (.A1(net3286),
    .A2(net3270),
    .B(net3269),
    .Y(_06098_));
 INVx1_ASAP7_75t_R _12220_ (.A(_06084_),
    .Y(_06099_));
 XOR2x2_ASAP7_75t_R _12221_ (.A(net3268),
    .B(_06098_),
    .Y(_06100_));
 AOI21x1_ASAP7_75t_R _12222_ (.A1(_06088_),
    .A2(_06097_),
    .B(_06058_),
    .Y(_06101_));
 XOR2x2_ASAP7_75t_R _12223_ (.A(_06089_),
    .B(net4246),
    .Y(_06102_));
 AO21x1_ASAP7_75t_R _12224_ (.A1(_06076_),
    .A2(_06068_),
    .B(_06089_),
    .Y(_06103_));
 OAI21x1_ASAP7_75t_R _12225_ (.A1(net3303),
    .A2(_06102_),
    .B(_06103_),
    .Y(_06104_));
 XNOR2x2_ASAP7_75t_R _12226_ (.A(net3284),
    .B(_06104_),
    .Y(_06105_));
 NAND2x1p5_ASAP7_75t_R _12227_ (.A(_06101_),
    .B(net3283),
    .Y(_06106_));
 OAI21x1_ASAP7_75t_R _12228_ (.A1(net3251),
    .A2(_06105_),
    .B(_06106_),
    .Y(_06107_));
 NOR2x1p5_ASAP7_75t_R _12229_ (.A(_06100_),
    .B(_06107_),
    .Y(_06108_));
 OR3x1_ASAP7_75t_R _12230_ (.A(net4504),
    .B(net4506),
    .C(_05574_),
    .Y(_06109_));
 XNOR2x2_ASAP7_75t_R _12231_ (.A(net4497),
    .B(_06109_),
    .Y(_06110_));
 NAND2x1p5_ASAP7_75t_R _12232_ (.A(_06101_),
    .B(net4244),
    .Y(_06111_));
 AOI211x1_ASAP7_75t_R _12233_ (.A1(net3302),
    .A2(_06091_),
    .B(net3368),
    .C(net4180),
    .Y(_06112_));
 XOR2x2_ASAP7_75t_R _12234_ (.A(_06055_),
    .B(net3359),
    .Y(_06113_));
 NAND2x1_ASAP7_75t_R _12235_ (.A(_06113_),
    .B(_06099_),
    .Y(_06114_));
 INVx1_ASAP7_75t_R _12236_ (.A(_06058_),
    .Y(_06115_));
 OAI21x1_ASAP7_75t_R _12237_ (.A1(_06112_),
    .A2(_06114_),
    .B(_06115_),
    .Y(_06116_));
 NAND2x1_ASAP7_75t_R _12238_ (.A(net4181),
    .B(_06116_),
    .Y(_06117_));
 NAND2x1_ASAP7_75t_R _12239_ (.A(net3323),
    .B(net3302),
    .Y(_06118_));
 INVx1_ASAP7_75t_R _12240_ (.A(_06118_),
    .Y(_06119_));
 AOI21x1_ASAP7_75t_R _12241_ (.A1(_06111_),
    .A2(_06117_),
    .B(_06119_),
    .Y(_06120_));
 NAND2x1p5_ASAP7_75t_R _12242_ (.A(_06110_),
    .B(_06120_),
    .Y(_06121_));
 AO21x1_ASAP7_75t_R _12243_ (.A1(_06120_),
    .A2(net4301),
    .B(net3227),
    .Y(_06122_));
 NOR2x1_ASAP7_75t_R _12244_ (.A(net3285),
    .B(net3282),
    .Y(_06123_));
 AO21x1_ASAP7_75t_R _12245_ (.A1(_06123_),
    .A2(net3286),
    .B(_06113_),
    .Y(_06124_));
 NAND2x1_ASAP7_75t_R _12246_ (.A(net3269),
    .B(net3270),
    .Y(_06125_));
 AND2x2_ASAP7_75t_R _12247_ (.A(_06124_),
    .B(_06125_),
    .Y(_06126_));
 INVx1_ASAP7_75t_R _12248_ (.A(_06126_),
    .Y(_06127_));
 OA21x2_ASAP7_75t_R _12249_ (.A1(_06122_),
    .A2(net3225),
    .B(net5619),
    .Y(_06128_));
 AOI21x1_ASAP7_75t_R _12250_ (.A1(net3213),
    .A2(net3195),
    .B(_06128_),
    .Y(_06129_));
 AOI21x1_ASAP7_75t_R _12251_ (.A1(_06108_),
    .A2(_06121_),
    .B(_06126_),
    .Y(_06130_));
 NOR2x1_ASAP7_75t_R _12252_ (.A(_06101_),
    .B(_06105_),
    .Y(_06131_));
 INVx1_ASAP7_75t_R _12253_ (.A(_06106_),
    .Y(_06132_));
 NOR2x1_ASAP7_75t_R _12254_ (.A(_06131_),
    .B(_06132_),
    .Y(_06133_));
 XOR2x2_ASAP7_75t_R _12255_ (.A(net3196),
    .B(net3212),
    .Y(_06134_));
 NOR2x1_ASAP7_75t_R _12256_ (.A(net3212),
    .B(net3238),
    .Y(_06135_));
 INVx1_ASAP7_75t_R _12257_ (.A(_06135_),
    .Y(_06136_));
 OAI21x1_ASAP7_75t_R _12258_ (.A1(net3185),
    .A2(_06134_),
    .B(_06136_),
    .Y(_06137_));
 XOR2x2_ASAP7_75t_R _12259_ (.A(_06118_),
    .B(net4181),
    .Y(_06138_));
 NAND2x1_ASAP7_75t_R _12260_ (.A(net3281),
    .B(net3251),
    .Y(_06139_));
 OA21x2_ASAP7_75t_R _12261_ (.A1(net3251),
    .A2(_06138_),
    .B(_06139_),
    .Y(_06140_));
 INVx1_ASAP7_75t_R _12262_ (.A(_06140_),
    .Y(_06141_));
 NAND2x1_ASAP7_75t_R _12263_ (.A(_06130_),
    .B(_06141_),
    .Y(_06142_));
 NOR2x1_ASAP7_75t_R _12264_ (.A(_06101_),
    .B(net4244),
    .Y(_06143_));
 NOR2x1_ASAP7_75t_R _12265_ (.A(net4181),
    .B(_06116_),
    .Y(_06144_));
 OAI21x1_ASAP7_75t_R _12266_ (.A1(net3237),
    .A2(net3224),
    .B(net4301),
    .Y(_06145_));
 XOR2x2_ASAP7_75t_R _12267_ (.A(_06140_),
    .B(_06145_),
    .Y(_06146_));
 INVx1_ASAP7_75t_R _12268_ (.A(_06100_),
    .Y(_06147_));
 NAND2x1_ASAP7_75t_R _12269_ (.A(_06147_),
    .B(_06133_),
    .Y(_06148_));
 INVx1_ASAP7_75t_R _12270_ (.A(_06110_),
    .Y(_06149_));
 OAI21x1_ASAP7_75t_R _12271_ (.A1(_06144_),
    .A2(_06143_),
    .B(net3281),
    .Y(_06150_));
 NOR2x1_ASAP7_75t_R _12272_ (.A(_06149_),
    .B(_06150_),
    .Y(_06151_));
 OAI21x1_ASAP7_75t_R _12273_ (.A1(_06148_),
    .A2(_06151_),
    .B(_06127_),
    .Y(_06152_));
 NAND2x1_ASAP7_75t_R _12274_ (.A(_06146_),
    .B(_06152_),
    .Y(_06153_));
 NAND2x1p5_ASAP7_75t_R _12275_ (.A(_06153_),
    .B(_06142_),
    .Y(_06154_));
 NOR2x2_ASAP7_75t_R _12276_ (.A(_06137_),
    .B(_06154_),
    .Y(_06155_));
 OR3x1_ASAP7_75t_R _12277_ (.A(net4504),
    .B(net4506),
    .C(_05655_),
    .Y(_06156_));
 XNOR2x2_ASAP7_75t_R _12278_ (.A(net4539),
    .B(_06156_),
    .Y(_06157_));
 NAND2x1_ASAP7_75t_R _12279_ (.A(net4300),
    .B(_06130_),
    .Y(_06158_));
 NAND2x1_ASAP7_75t_R _12280_ (.A(_06152_),
    .B(net4243),
    .Y(_06159_));
 NAND2x1_ASAP7_75t_R _12281_ (.A(net3239),
    .B(net3226),
    .Y(_06160_));
 INVx1_ASAP7_75t_R _12282_ (.A(net3207),
    .Y(_06161_));
 AOI21x1_ASAP7_75t_R _12283_ (.A1(_06158_),
    .A2(_06159_),
    .B(_06161_),
    .Y(_06162_));
 NAND2x1_ASAP7_75t_R _12284_ (.A(_06162_),
    .B(_06157_),
    .Y(_06163_));
 OAI21x1_ASAP7_75t_R _12285_ (.A1(net3177),
    .A2(_06155_),
    .B(net3146),
    .Y(_06164_));
 XOR2x2_ASAP7_75t_R _12286_ (.A(_06164_),
    .B(net3162),
    .Y(_06165_));
 XOR2x2_ASAP7_75t_R _12287_ (.A(_06160_),
    .B(net4243),
    .Y(_06166_));
 NAND2x1_ASAP7_75t_R _12288_ (.A(net3208),
    .B(net3185),
    .Y(_06167_));
 OAI21x1_ASAP7_75t_R _12289_ (.A1(net3185),
    .A2(_06166_),
    .B(_06167_),
    .Y(_06168_));
 INVx1_ASAP7_75t_R _12290_ (.A(net3161),
    .Y(_06169_));
 INVx1_ASAP7_75t_R _12291_ (.A(net3210),
    .Y(_06170_));
 AOI21x1_ASAP7_75t_R _12292_ (.A1(_06170_),
    .A2(_06152_),
    .B(net3211),
    .Y(_06171_));
 NOR2x1_ASAP7_75t_R _12293_ (.A(net3195),
    .B(net3185),
    .Y(_06172_));
 XOR2x2_ASAP7_75t_R _12294_ (.A(net3197),
    .B(net3227),
    .Y(_06173_));
 AOI21x1_ASAP7_75t_R _12295_ (.A1(net5605),
    .A2(_06173_),
    .B(net3194),
    .Y(_06174_));
 OAI21x1_ASAP7_75t_R _12296_ (.A1(_06171_),
    .A2(_06172_),
    .B(_06174_),
    .Y(_06175_));
 INVx1_ASAP7_75t_R _12297_ (.A(_06157_),
    .Y(_06176_));
 AOI211x1_ASAP7_75t_R _12298_ (.A1(net3213),
    .A2(net3209),
    .B(net3238),
    .C(net4243),
    .Y(_06177_));
 NAND2x1_ASAP7_75t_R _12299_ (.A(net3213),
    .B(net3195),
    .Y(_06178_));
 AOI21x1_ASAP7_75t_R _12300_ (.A1(net3225),
    .A2(_06178_),
    .B(net4300),
    .Y(_06179_));
 OAI21x1_ASAP7_75t_R _12301_ (.A1(_06177_),
    .A2(_06179_),
    .B(net3207),
    .Y(_06180_));
 NOR2x1_ASAP7_75t_R _12302_ (.A(_06176_),
    .B(_06180_),
    .Y(_06181_));
 INVx1_ASAP7_75t_R _12303_ (.A(_06129_),
    .Y(_06182_));
 OAI21x1_ASAP7_75t_R _12304_ (.A1(_06175_),
    .A2(_06181_),
    .B(_06182_),
    .Y(_06183_));
 NOR2x1_ASAP7_75t_R _12305_ (.A(_06169_),
    .B(_06183_),
    .Y(_06184_));
 OAI21x1_ASAP7_75t_R _12306_ (.A1(_06177_),
    .A2(_06179_),
    .B(_06157_),
    .Y(_06185_));
 XNOR2x2_ASAP7_75t_R _12307_ (.A(_06168_),
    .B(_06185_),
    .Y(_06186_));
 INVx1_ASAP7_75t_R _12308_ (.A(_06186_),
    .Y(_06187_));
 AOI21x1_ASAP7_75t_R _12309_ (.A1(_06155_),
    .A2(_06163_),
    .B(_06129_),
    .Y(_06188_));
 NOR2x1_ASAP7_75t_R _12310_ (.A(_06188_),
    .B(_06187_),
    .Y(_06189_));
 NOR2x1_ASAP7_75t_R _12311_ (.A(_06189_),
    .B(_06184_),
    .Y(_06190_));
 NAND2x1_ASAP7_75t_R _12312_ (.A(_06190_),
    .B(_06165_),
    .Y(_06191_));
 AOI211x1_ASAP7_75t_R _12313_ (.A1(net5634),
    .A2(net3160),
    .B(net3177),
    .C(net4241),
    .Y(_06192_));
 OAI21x1_ASAP7_75t_R _12314_ (.A1(net4241),
    .A2(net3160),
    .B(net5634),
    .Y(_06193_));
 AOI21x1_ASAP7_75t_R _12315_ (.A1(_06182_),
    .A2(_06193_),
    .B(net4299),
    .Y(_06194_));
 NAND2x1_ASAP7_75t_R _12316_ (.A(net3175),
    .B(net3174),
    .Y(_06195_));
 OAI21x1_ASAP7_75t_R _12317_ (.A1(_06194_),
    .A2(_06192_),
    .B(_06195_),
    .Y(_06196_));
 NOR2x1p5_ASAP7_75t_R _12318_ (.A(_05491_),
    .B(_06196_),
    .Y(_06197_));
 AO21x1_ASAP7_75t_R _12319_ (.A1(_06162_),
    .A2(_06157_),
    .B(net3162),
    .Y(_06198_));
 OA21x2_ASAP7_75t_R _12320_ (.A1(_06198_),
    .A2(net3159),
    .B(net3176),
    .Y(_06199_));
 AOI21x1_ASAP7_75t_R _12321_ (.A1(net3147),
    .A2(net3148),
    .B(_06199_),
    .Y(_06200_));
 INVx1_ASAP7_75t_R _12322_ (.A(_06200_),
    .Y(_06201_));
 OAI21x1_ASAP7_75t_R _12323_ (.A1(_06197_),
    .A2(_06191_),
    .B(_06201_),
    .Y(_06202_));
 NAND2x1_ASAP7_75t_R _12324_ (.A(net4253),
    .B(_06202_),
    .Y(_06203_));
 XNOR2x2_ASAP7_75t_R _12325_ (.A(net3162),
    .B(_06164_),
    .Y(_06204_));
 NAND2x1_ASAP7_75t_R _12326_ (.A(net3145),
    .B(_06183_),
    .Y(_06205_));
 NAND2x1_ASAP7_75t_R _12327_ (.A(net3161),
    .B(_06188_),
    .Y(_06206_));
 NAND2x1_ASAP7_75t_R _12328_ (.A(_06205_),
    .B(_06206_),
    .Y(_06207_));
 NOR2x1p5_ASAP7_75t_R _12329_ (.A(_06204_),
    .B(_06207_),
    .Y(_06208_));
 NAND2x1_ASAP7_75t_R _12330_ (.A(net4242),
    .B(net3134),
    .Y(_06209_));
 NAND2x1_ASAP7_75t_R _12331_ (.A(net4299),
    .B(net3133),
    .Y(_06210_));
 INVx1_ASAP7_75t_R _12332_ (.A(net3158),
    .Y(_06211_));
 AOI21x1_ASAP7_75t_R _12333_ (.A1(_06209_),
    .A2(_06210_),
    .B(_06211_),
    .Y(_06212_));
 NAND2x1_ASAP7_75t_R _12334_ (.A(net4308),
    .B(_06212_),
    .Y(_06213_));
 AOI21x1_ASAP7_75t_R _12335_ (.A1(_06208_),
    .A2(_06213_),
    .B(net3122),
    .Y(_06214_));
 NAND2x1_ASAP7_75t_R _12336_ (.A(net4308),
    .B(_06214_),
    .Y(_06215_));
 NAND2x1_ASAP7_75t_R _12337_ (.A(_06215_),
    .B(_06203_),
    .Y(_06216_));
 INVx1_ASAP7_75t_R _12338_ (.A(_06216_),
    .Y(_06217_));
 NOR2x1_ASAP7_75t_R _12339_ (.A(_05478_),
    .B(_06217_),
    .Y(_06218_));
 INVx1_ASAP7_75t_R _12340_ (.A(_06218_),
    .Y(_06219_));
 NAND2x1_ASAP7_75t_R _12341_ (.A(net4308),
    .B(net3088),
    .Y(_06220_));
 NAND2x1_ASAP7_75t_R _12342_ (.A(net3120),
    .B(net3119),
    .Y(_06221_));
 XOR2x2_ASAP7_75t_R _12343_ (.A(_06220_),
    .B(net3109),
    .Y(_06222_));
 OAI21x1_ASAP7_75t_R _12344_ (.A1(net3122),
    .A2(_06208_),
    .B(_06213_),
    .Y(_06223_));
 XOR2x2_ASAP7_75t_R _12345_ (.A(_06223_),
    .B(net3113),
    .Y(_06224_));
 XOR2x2_ASAP7_75t_R _12346_ (.A(_06195_),
    .B(net4242),
    .Y(_06225_));
 NAND2x1_ASAP7_75t_R _12347_ (.A(net3158),
    .B(net3133),
    .Y(_06226_));
 OAI21x1_ASAP7_75t_R _12348_ (.A1(net3133),
    .A2(_06225_),
    .B(_06226_),
    .Y(_06227_));
 INVx1_ASAP7_75t_R _12349_ (.A(net3108),
    .Y(_06228_));
 OAI21x1_ASAP7_75t_R _12350_ (.A1(net3132),
    .A2(net3123),
    .B(net4308),
    .Y(_06229_));
 XNOR2x2_ASAP7_75t_R _12351_ (.A(_06227_),
    .B(_06229_),
    .Y(_06230_));
 NAND2x1_ASAP7_75t_R _12352_ (.A(_06230_),
    .B(_06202_),
    .Y(_06231_));
 OAI21x1_ASAP7_75t_R _12353_ (.A1(_06228_),
    .A2(net3089),
    .B(_06231_),
    .Y(_06232_));
 NOR2x1_ASAP7_75t_R _12354_ (.A(_06232_),
    .B(_06224_),
    .Y(_06233_));
 NOR2x1_ASAP7_75t_R _12355_ (.A(net3110),
    .B(net3099),
    .Y(_06234_));
 NAND2x1_ASAP7_75t_R _12356_ (.A(_06234_),
    .B(_06202_),
    .Y(_06235_));
 OAI21x1_ASAP7_75t_R _12357_ (.A1(net4253),
    .A2(net3112),
    .B(_06208_),
    .Y(_06236_));
 INVx1_ASAP7_75t_R _12358_ (.A(_06236_),
    .Y(_06237_));
 AOI21x1_ASAP7_75t_R _12359_ (.A1(_06235_),
    .A2(net3121),
    .B(_06237_),
    .Y(_06238_));
 AOI21x1_ASAP7_75t_R _12360_ (.A1(_06222_),
    .A2(net3043),
    .B(net3059),
    .Y(_06239_));
 OAI21x1_ASAP7_75t_R _12361_ (.A1(_06219_),
    .A2(_06239_),
    .B(_06222_),
    .Y(_06240_));
 INVx2_ASAP7_75t_R _12362_ (.A(_06238_),
    .Y(_06241_));
 INVx1_ASAP7_75t_R _12363_ (.A(_06221_),
    .Y(_06242_));
 AOI21x1_ASAP7_75t_R _12364_ (.A1(_06203_),
    .A2(_06215_),
    .B(_06242_),
    .Y(_06243_));
 NAND2x1_ASAP7_75t_R _12365_ (.A(_05477_),
    .B(_06243_),
    .Y(_06244_));
 NOR2x1_ASAP7_75t_R _12366_ (.A(_06241_),
    .B(net3041),
    .Y(_06245_));
 INVx1_ASAP7_75t_R _12367_ (.A(_06245_),
    .Y(_06246_));
 AOI211x1_ASAP7_75t_R _12368_ (.A1(net3098),
    .A2(net3112),
    .B(net3122),
    .C(net4253),
    .Y(_06247_));
 AOI21x1_ASAP7_75t_R _12369_ (.A1(net3111),
    .A2(net3085),
    .B(net4308),
    .Y(_06248_));
 OAI21x1_ASAP7_75t_R _12370_ (.A1(_06247_),
    .A2(_06248_),
    .B(net3109),
    .Y(_06249_));
 NOR2x1_ASAP7_75t_R _12371_ (.A(_05478_),
    .B(_06249_),
    .Y(_06250_));
 OAI21x1_ASAP7_75t_R _12372_ (.A1(_06241_),
    .A2(_06250_),
    .B(net3060),
    .Y(_06251_));
 NOR2x1_ASAP7_75t_R _12373_ (.A(net3075),
    .B(_06238_),
    .Y(_06252_));
 AOI21x1_ASAP7_75t_R _12374_ (.A1(net4309),
    .A2(net3057),
    .B(net5621),
    .Y(_06253_));
 OAI21x1_ASAP7_75t_R _12375_ (.A1(net3058),
    .A2(_06252_),
    .B(_06253_),
    .Y(_06254_));
 NAND2x1_ASAP7_75t_R _12376_ (.A(_06251_),
    .B(_06254_),
    .Y(_06255_));
 AOI21x1_ASAP7_75t_R _12377_ (.A1(_06240_),
    .A2(_06246_),
    .B(_06255_),
    .Y(_06256_));
 AOI211x1_ASAP7_75t_R _12378_ (.A1(_06233_),
    .A2(_06249_),
    .B(net3059),
    .C(net4254),
    .Y(_06257_));
 AOI21x1_ASAP7_75t_R _12379_ (.A1(_06244_),
    .A2(_06233_),
    .B(_06238_),
    .Y(_06258_));
 NOR2x1_ASAP7_75t_R _12380_ (.A(net4310),
    .B(_06258_),
    .Y(_06259_));
 OAI21x1_ASAP7_75t_R _12381_ (.A1(_06257_),
    .A2(_06259_),
    .B(net3061),
    .Y(_06260_));
 XOR2x2_ASAP7_75t_R _12382_ (.A(net3086),
    .B(net3110),
    .Y(_06261_));
 XOR2x2_ASAP7_75t_R _12383_ (.A(_06254_),
    .B(net3074),
    .Y(_06262_));
 INVx3_ASAP7_75t_R _12384_ (.A(_06262_),
    .Y(_06263_));
 BUFx3_ASAP7_75t_R place2938 (.A(_06314_),
    .Y(net2938));
 NOR2x1_ASAP7_75t_R _12386_ (.A(net4502),
    .B(net4400),
    .Y(_06265_));
 XOR2x2_ASAP7_75t_R _12387_ (.A(_06265_),
    .B(net4508),
    .Y(_06266_));
 INVx1_ASAP7_75t_R _12388_ (.A(_06266_),
    .Y(_06267_));
 AOI211x1_ASAP7_75t_R _12389_ (.A1(_06260_),
    .A2(_06256_),
    .B(net4240),
    .C(_06263_),
    .Y(_06268_));
 OAI21x1_ASAP7_75t_R _12390_ (.A1(_06260_),
    .A2(_06267_),
    .B(_06256_),
    .Y(_06269_));
 AOI21x1_ASAP7_75t_R _12391_ (.A1(net3018),
    .A2(net5615),
    .B(net4298),
    .Y(_06270_));
 NOR2x1_ASAP7_75t_R _12392_ (.A(net4507),
    .B(net4400),
    .Y(_06271_));
 XOR2x2_ASAP7_75t_R _12393_ (.A(_06271_),
    .B(net4604),
    .Y(_06272_));
 OAI21x1_ASAP7_75t_R _12394_ (.A1(net2986),
    .A2(_06270_),
    .B(net4296),
    .Y(_06273_));
 NOR2x1_ASAP7_75t_R _12395_ (.A(_06228_),
    .B(net3089),
    .Y(_06274_));
 INVx1_ASAP7_75t_R _12396_ (.A(_06230_),
    .Y(_06275_));
 NOR2x1_ASAP7_75t_R _12397_ (.A(_06275_),
    .B(net3087),
    .Y(_06276_));
 NOR2x1_ASAP7_75t_R _12398_ (.A(_06274_),
    .B(_06276_),
    .Y(_06277_));
 NAND2x1_ASAP7_75t_R _12399_ (.A(_06261_),
    .B(_06277_),
    .Y(_06278_));
 OAI21x1_ASAP7_75t_R _12400_ (.A1(_06278_),
    .A2(_06250_),
    .B(_06241_),
    .Y(_06279_));
 NAND2x1_ASAP7_75t_R _12401_ (.A(net4255),
    .B(_06279_),
    .Y(_06280_));
 NAND2x1_ASAP7_75t_R _12402_ (.A(net4310),
    .B(net5602),
    .Y(_06281_));
 NAND2x1_ASAP7_75t_R _12403_ (.A(_06280_),
    .B(_06281_),
    .Y(_06282_));
 INVx1_ASAP7_75t_R _12404_ (.A(net3010),
    .Y(_06283_));
 NAND2x1_ASAP7_75t_R _12405_ (.A(net3018),
    .B(_06269_),
    .Y(_06284_));
 INVx1_ASAP7_75t_R _12406_ (.A(_06269_),
    .Y(_06285_));
 XOR2x2_ASAP7_75t_R _12407_ (.A(_06282_),
    .B(net4298),
    .Y(_06286_));
 OAI21x1_ASAP7_75t_R _12408_ (.A1(net3011),
    .A2(net2974),
    .B(_06286_),
    .Y(_06287_));
 OAI21x1_ASAP7_75t_R _12409_ (.A1(_06283_),
    .A2(net2975),
    .B(_06287_),
    .Y(_06288_));
 XNOR2x2_ASAP7_75t_R _12410_ (.A(_06273_),
    .B(_06288_),
    .Y(_06289_));
 OAI21x1_ASAP7_75t_R _12411_ (.A1(_06257_),
    .A2(_06259_),
    .B(_06266_),
    .Y(_06290_));
 NOR2x1_ASAP7_75t_R _12412_ (.A(net3044),
    .B(_06279_),
    .Y(_06291_));
 XOR2x2_ASAP7_75t_R _12413_ (.A(net5924),
    .B(_05478_),
    .Y(_06292_));
 NOR2x1_ASAP7_75t_R _12414_ (.A(_06292_),
    .B(net5626),
    .Y(_06293_));
 NOR2x1_ASAP7_75t_R _12415_ (.A(_06291_),
    .B(_06293_),
    .Y(_06294_));
 XOR2x2_ASAP7_75t_R _12416_ (.A(_06294_),
    .B(_06290_),
    .Y(_06295_));
 AOI211x1_ASAP7_75t_R _12417_ (.A1(_06256_),
    .A2(_06290_),
    .B(_06263_),
    .C(net3009),
    .Y(_06296_));
 AOI21x1_ASAP7_75t_R _12418_ (.A1(_06284_),
    .A2(_06295_),
    .B(_06296_),
    .Y(_06297_));
 XOR2x2_ASAP7_75t_R _12419_ (.A(_06220_),
    .B(net3097),
    .Y(_06298_));
 OAI21x1_ASAP7_75t_R _12420_ (.A1(_06298_),
    .A2(_06278_),
    .B(net3042),
    .Y(_06299_));
 AOI21x1_ASAP7_75t_R _12421_ (.A1(_06218_),
    .A2(_06299_),
    .B(_06298_),
    .Y(_06300_));
 AOI21x1_ASAP7_75t_R _12422_ (.A1(net3058),
    .A2(net3041),
    .B(net3055),
    .Y(_06301_));
 OAI21x1_ASAP7_75t_R _12423_ (.A1(net4254),
    .A2(net3056),
    .B(net3055),
    .Y(_06302_));
 AOI21x1_ASAP7_75t_R _12424_ (.A1(net3042),
    .A2(net3075),
    .B(_06302_),
    .Y(_06303_));
 NOR2x1_ASAP7_75t_R _12425_ (.A(_06301_),
    .B(_06303_),
    .Y(_06304_));
 OAI21x1_ASAP7_75t_R _12426_ (.A1(_06300_),
    .A2(net3031),
    .B(_06304_),
    .Y(_06305_));
 AOI21x1_ASAP7_75t_R _12427_ (.A1(_06280_),
    .A2(_06281_),
    .B(net3044),
    .Y(_06306_));
 AOI22x1_ASAP7_75t_R _12428_ (.A1(_06305_),
    .A2(_06262_),
    .B1(net4298),
    .B2(_06306_),
    .Y(_06307_));
 NOR2x1_ASAP7_75t_R _12429_ (.A(net3031),
    .B(_06300_),
    .Y(_06308_));
 INVx1_ASAP7_75t_R _12430_ (.A(_06308_),
    .Y(_06309_));
 XOR2x2_ASAP7_75t_R _12431_ (.A(_06307_),
    .B(net2997),
    .Y(_06310_));
 NAND2x1_ASAP7_75t_R _12432_ (.A(_06297_),
    .B(_06310_),
    .Y(_06311_));
 INVx1_ASAP7_75t_R _12433_ (.A(_06272_),
    .Y(_06312_));
 OAI21x1_ASAP7_75t_R _12434_ (.A1(_06270_),
    .A2(_06268_),
    .B(net3010),
    .Y(_06313_));
 NOR2x1p5_ASAP7_75t_R _12435_ (.A(_06312_),
    .B(_06313_),
    .Y(_06314_));
 OA21x2_ASAP7_75t_R _12436_ (.A1(net5597),
    .A2(net4240),
    .B(_06309_),
    .Y(_06315_));
 NOR2x1_ASAP7_75t_R _12437_ (.A(net3017),
    .B(_06315_),
    .Y(_06316_));
 AO21x1_ASAP7_75t_R _12438_ (.A1(_06315_),
    .A2(net3019),
    .B(_06316_),
    .Y(_06317_));
 OAI21x1_ASAP7_75t_R _12439_ (.A1(_06314_),
    .A2(_06311_),
    .B(net2957),
    .Y(_06318_));
 NAND2x1_ASAP7_75t_R _12440_ (.A(_06318_),
    .B(_06289_),
    .Y(_06319_));
 XOR2x2_ASAP7_75t_R _12441_ (.A(_06307_),
    .B(net3008),
    .Y(_06320_));
 INVx1_ASAP7_75t_R _12442_ (.A(_06296_),
    .Y(_06321_));
 OAI21x1_ASAP7_75t_R _12443_ (.A1(net3011),
    .A2(_06285_),
    .B(_06295_),
    .Y(_06322_));
 NAND2x1_ASAP7_75t_R _12444_ (.A(_06322_),
    .B(_06321_),
    .Y(_06323_));
 NOR2x1_ASAP7_75t_R _12445_ (.A(_06320_),
    .B(_06323_),
    .Y(_06324_));
 NOR2x1_ASAP7_75t_R _12446_ (.A(net5597),
    .B(_06305_),
    .Y(_06325_));
 OAI21x1_ASAP7_75t_R _12447_ (.A1(_06306_),
    .A2(_06305_),
    .B(_06262_),
    .Y(_06326_));
 OAI21x1_ASAP7_75t_R _12448_ (.A1(_06326_),
    .A2(_06325_),
    .B(net4240),
    .Y(_06327_));
 INVx1_ASAP7_75t_R _12449_ (.A(_06268_),
    .Y(_06328_));
 AOI21x1_ASAP7_75t_R _12450_ (.A1(_06327_),
    .A2(_06328_),
    .B(_06283_),
    .Y(_06329_));
 NAND2x1_ASAP7_75t_R _12451_ (.A(net4296),
    .B(_06329_),
    .Y(_06330_));
 INVx2_ASAP7_75t_R _12452_ (.A(_06317_),
    .Y(_06331_));
 AOI21x1_ASAP7_75t_R _12453_ (.A1(_06330_),
    .A2(_06324_),
    .B(_06331_),
    .Y(_06332_));
 NAND2x1_ASAP7_75t_R _12454_ (.A(_06332_),
    .B(net2940),
    .Y(_06333_));
 NAND2x1p5_ASAP7_75t_R _12455_ (.A(_06319_),
    .B(_06333_),
    .Y(_06334_));
 NOR2x1_ASAP7_75t_R _12456_ (.A(net2937),
    .B(net2938),
    .Y(_06335_));
 NAND2x1_ASAP7_75t_R _12457_ (.A(_06335_),
    .B(_06318_),
    .Y(_06336_));
 NOR2x1_ASAP7_75t_R _12458_ (.A(net2939),
    .B(net2938),
    .Y(_06337_));
 AOI21x1_ASAP7_75t_R _12459_ (.A1(net2985),
    .A2(_06336_),
    .B(_06337_),
    .Y(_06338_));
 OAI21x1_ASAP7_75t_R _12460_ (.A1(_06331_),
    .A2(_06324_),
    .B(_06330_),
    .Y(_06339_));
 XOR2x2_ASAP7_75t_R _12461_ (.A(_06339_),
    .B(net2958),
    .Y(_06340_));
 NOR2x2_ASAP7_75t_R _12462_ (.A(_06334_),
    .B(_06340_),
    .Y(_06341_));
 NOR2x1_ASAP7_75t_R _12463_ (.A(net4547),
    .B(net4400),
    .Y(_06342_));
 XOR2x2_ASAP7_75t_R _12464_ (.A(_06342_),
    .B(net4605),
    .Y(_06343_));
 NAND2x1_ASAP7_75t_R _12465_ (.A(net4239),
    .B(_06318_),
    .Y(_06344_));
 NAND2x1_ASAP7_75t_R _12466_ (.A(net4297),
    .B(_06332_),
    .Y(_06345_));
 NAND2x1_ASAP7_75t_R _12467_ (.A(net2984),
    .B(net2973),
    .Y(_06346_));
 INVx1_ASAP7_75t_R _12468_ (.A(_06346_),
    .Y(_06347_));
 AOI21x1_ASAP7_75t_R _12469_ (.A1(_06344_),
    .A2(_06345_),
    .B(_06347_),
    .Y(_06348_));
 NAND2x1_ASAP7_75t_R _12470_ (.A(_06343_),
    .B(_06348_),
    .Y(_06349_));
 OAI21x1_ASAP7_75t_R _12471_ (.A1(_06338_),
    .A2(_06341_),
    .B(_06349_),
    .Y(_06350_));
 NOR2x1_ASAP7_75t_R _12472_ (.A(net2882),
    .B(_06350_),
    .Y(_06351_));
 XOR2x2_ASAP7_75t_R _12473_ (.A(_06351_),
    .B(net2897),
    .Y(_06352_));
 INVx2_ASAP7_75t_R _12474_ (.A(_06352_),
    .Y(_06353_));
 XOR2x2_ASAP7_75t_R _12475_ (.A(net2927),
    .B(net4239),
    .Y(_06354_));
 INVx1_ASAP7_75t_R _12476_ (.A(net2917),
    .Y(_06355_));
 INVx1_ASAP7_75t_R _12477_ (.A(net2881),
    .Y(_06356_));
 XOR2x2_ASAP7_75t_R _12478_ (.A(_06339_),
    .B(net2937),
    .Y(_06357_));
 INVx1_ASAP7_75t_R _12479_ (.A(net2940),
    .Y(_06358_));
 NOR2x1_ASAP7_75t_R _12480_ (.A(_06358_),
    .B(net2927),
    .Y(_06359_));
 XOR2x2_ASAP7_75t_R _12481_ (.A(net2940),
    .B(net2959),
    .Y(_06360_));
 NOR2x1_ASAP7_75t_R _12482_ (.A(_06360_),
    .B(net2918),
    .Y(_06361_));
 NOR2x1_ASAP7_75t_R _12483_ (.A(_06359_),
    .B(_06361_),
    .Y(_06362_));
 NAND2x1_ASAP7_75t_R _12484_ (.A(_06357_),
    .B(_06362_),
    .Y(_06363_));
 NOR2x1_ASAP7_75t_R _12485_ (.A(net2865),
    .B(_06363_),
    .Y(_06364_));
 INVx1_ASAP7_75t_R _12486_ (.A(_06338_),
    .Y(_06365_));
 OAI21x1_ASAP7_75t_R _12487_ (.A1(net2881),
    .A2(_06363_),
    .B(_06365_),
    .Y(_06366_));
 INVx1_ASAP7_75t_R _12488_ (.A(_06343_),
    .Y(_06367_));
 OAI21x1_ASAP7_75t_R _12489_ (.A1(_06364_),
    .A2(_06366_),
    .B(net4238),
    .Y(_06368_));
 AOI211x1_ASAP7_75t_R _12490_ (.A1(net2867),
    .A2(_06356_),
    .B(net2898),
    .C(net4238),
    .Y(_06369_));
 INVx1_ASAP7_75t_R _12491_ (.A(_06369_),
    .Y(_06370_));
 NOR2x1_ASAP7_75t_R _12492_ (.A(net4548),
    .B(net4400),
    .Y(_06371_));
 XOR2x2_ASAP7_75t_R _12493_ (.A(_06371_),
    .B(net4663),
    .Y(_06372_));
 INVx1_ASAP7_75t_R _12494_ (.A(_06372_),
    .Y(_06373_));
 AOI21x1_ASAP7_75t_R _12495_ (.A1(_06370_),
    .A2(_06368_),
    .B(_06373_),
    .Y(_06374_));
 AND3x2_ASAP7_75t_R _12496_ (.A(_06353_),
    .B(net2896),
    .C(net2824),
    .Y(_06375_));
 XOR2x2_ASAP7_75t_R _12497_ (.A(_06350_),
    .B(net2880),
    .Y(_06376_));
 XOR2x2_ASAP7_75t_R _12498_ (.A(_06346_),
    .B(net4297),
    .Y(_06377_));
 NAND2x1_ASAP7_75t_R _12499_ (.A(_06377_),
    .B(net2927),
    .Y(_06378_));
 OAI21x1_ASAP7_75t_R _12500_ (.A1(net2936),
    .A2(net2927),
    .B(_06378_),
    .Y(_06379_));
 INVx1_ASAP7_75t_R _12501_ (.A(_06379_),
    .Y(_06380_));
 NAND2x1_ASAP7_75t_R _12502_ (.A(_06380_),
    .B(net2867),
    .Y(_06381_));
 AO21x1_ASAP7_75t_R _12503_ (.A1(_06345_),
    .A2(_06344_),
    .B(_06367_),
    .Y(_06382_));
 AOI21x1_ASAP7_75t_R _12504_ (.A1(_06365_),
    .A2(_06381_),
    .B(net2878),
    .Y(_06383_));
 NOR2x1_ASAP7_75t_R _12505_ (.A(_06367_),
    .B(_06354_),
    .Y(_06384_));
 AND3x1_ASAP7_75t_R _12506_ (.A(_06384_),
    .B(net2956),
    .C(net2899),
    .Y(_06385_));
 INVx1_ASAP7_75t_R _12507_ (.A(_06385_),
    .Y(_06386_));
 OAI21x1_ASAP7_75t_R _12508_ (.A1(net2895),
    .A2(_06383_),
    .B(_06386_),
    .Y(_06387_));
 XOR2x2_ASAP7_75t_R _12509_ (.A(net2917),
    .B(net4295),
    .Y(_06388_));
 AOI21x1_ASAP7_75t_R _12510_ (.A1(net2868),
    .A2(net2866),
    .B(net2898),
    .Y(_06389_));
 NOR2x1_ASAP7_75t_R _12511_ (.A(_06388_),
    .B(_06389_),
    .Y(_06390_));
 AOI211x1_ASAP7_75t_R _12512_ (.A1(net2866),
    .A2(net2868),
    .B(net2917),
    .C(net2898),
    .Y(_06391_));
 NOR2x1_ASAP7_75t_R _12513_ (.A(_06390_),
    .B(_06391_),
    .Y(_06392_));
 NAND2x1_ASAP7_75t_R _12514_ (.A(_06387_),
    .B(_06392_),
    .Y(_06393_));
 OAI21x1_ASAP7_75t_R _12515_ (.A1(net2835),
    .A2(_06393_),
    .B(net2825),
    .Y(_06394_));
 INVx1_ASAP7_75t_R _12516_ (.A(_06392_),
    .Y(_06395_));
 AOI21x1_ASAP7_75t_R _12517_ (.A1(net2824),
    .A2(_06394_),
    .B(_06395_),
    .Y(_06396_));
 NOR2x1_ASAP7_75t_R _12518_ (.A(_06396_),
    .B(_06375_),
    .Y(_06397_));
 NOR2x1_ASAP7_75t_R _12519_ (.A(net4661),
    .B(net4400),
    .Y(_06398_));
 XOR2x2_ASAP7_75t_R _12520_ (.A(_06398_),
    .B(net4665),
    .Y(_06399_));
 NOR3x1_ASAP7_75t_R _12521_ (.A(_06379_),
    .B(net2882),
    .C(net2897),
    .Y(_06400_));
 OAI21x1_ASAP7_75t_R _12522_ (.A1(net2899),
    .A2(_06400_),
    .B(net2894),
    .Y(_06401_));
 AOI21x1_ASAP7_75t_R _12523_ (.A1(net2879),
    .A2(_06401_),
    .B(_06385_),
    .Y(_06402_));
 NOR2x1_ASAP7_75t_R _12524_ (.A(_06376_),
    .B(_06402_),
    .Y(_06403_));
 OA21x2_ASAP7_75t_R _12525_ (.A1(_06353_),
    .A2(_06403_),
    .B(net4237),
    .Y(_06404_));
 OAI21x1_ASAP7_75t_R _12526_ (.A1(net2936),
    .A2(_06382_),
    .B(net2867),
    .Y(_06405_));
 AOI21x1_ASAP7_75t_R _12527_ (.A1(_06365_),
    .A2(_06405_),
    .B(net4295),
    .Y(_06406_));
 OAI21x1_ASAP7_75t_R _12528_ (.A1(_06406_),
    .A2(_06369_),
    .B(_06355_),
    .Y(_06407_));
 AOI211x1_ASAP7_75t_R _12529_ (.A1(_06403_),
    .A2(_06407_),
    .B(_06353_),
    .C(net4237),
    .Y(_06408_));
 NOR2x1_ASAP7_75t_R _12530_ (.A(net2848),
    .B(net2834),
    .Y(_06409_));
 INVx1_ASAP7_75t_R _12531_ (.A(_06409_),
    .Y(_06410_));
 OAI21x1_ASAP7_75t_R _12532_ (.A1(_06408_),
    .A2(_06404_),
    .B(_06410_),
    .Y(_06411_));
 NOR2x1p5_ASAP7_75t_R _12533_ (.A(_06399_),
    .B(_06411_),
    .Y(_06412_));
 NOR2x1_ASAP7_75t_R _12534_ (.A(_06397_),
    .B(net2770),
    .Y(_06413_));
 INVx1_ASAP7_75t_R _12535_ (.A(_06397_),
    .Y(_06414_));
 NOR3x1_ASAP7_75t_R _12536_ (.A(_06414_),
    .B(net2784),
    .C(net4293),
    .Y(_06415_));
 NAND2x1_ASAP7_75t_R _12537_ (.A(_06374_),
    .B(net2896),
    .Y(_06416_));
 AOI21x1_ASAP7_75t_R _12538_ (.A1(_06353_),
    .A2(_06416_),
    .B(net2823),
    .Y(_06417_));
 OAI21x1_ASAP7_75t_R _12539_ (.A1(net4237),
    .A2(_06407_),
    .B(_06387_),
    .Y(_06418_));
 AOI21x1_ASAP7_75t_R _12540_ (.A1(net2835),
    .A2(net2825),
    .B(_06418_),
    .Y(_06419_));
 NOR2x1_ASAP7_75t_R _12541_ (.A(_06417_),
    .B(_06419_),
    .Y(_06420_));
 OAI21x1_ASAP7_75t_R _12542_ (.A1(_06375_),
    .A2(_06396_),
    .B(_06420_),
    .Y(_06421_));
 XOR2x2_ASAP7_75t_R _12543_ (.A(_06419_),
    .B(net2835),
    .Y(_06422_));
 OAI21x1_ASAP7_75t_R _12544_ (.A1(_06412_),
    .A2(_06421_),
    .B(_06422_),
    .Y(_06423_));
 OAI21x1_ASAP7_75t_R _12545_ (.A1(_06413_),
    .A2(_06415_),
    .B(net2758),
    .Y(_06424_));
 INVx1_ASAP7_75t_R _12546_ (.A(_06424_),
    .Y(_06425_));
 NOR2x2_ASAP7_75t_R _12547_ (.A(net2759),
    .B(net2758),
    .Y(_06426_));
 XOR2x2_ASAP7_75t_R _12548_ (.A(net2849),
    .B(net2882),
    .Y(_06427_));
 NAND2x1_ASAP7_75t_R _12549_ (.A(_06427_),
    .B(_06387_),
    .Y(_06428_));
 NOR2x1_ASAP7_75t_R _12550_ (.A(net4237),
    .B(_06407_),
    .Y(_06429_));
 OAI21x1_ASAP7_75t_R _12551_ (.A1(_06428_),
    .A2(_06429_),
    .B(net5664),
    .Y(_06430_));
 NOR2x1_ASAP7_75t_R _12552_ (.A(net4294),
    .B(net2822),
    .Y(_06431_));
 AND3x1_ASAP7_75t_R _12553_ (.A(net2836),
    .B(_06368_),
    .C(net4294),
    .Y(_06432_));
 OAI21x1_ASAP7_75t_R _12554_ (.A1(_06431_),
    .A2(_06432_),
    .B(_06430_),
    .Y(_06433_));
 OAI21x1_ASAP7_75t_R _12555_ (.A1(net2822),
    .A2(_06430_),
    .B(_06433_),
    .Y(_06434_));
 INVx1_ASAP7_75t_R _12556_ (.A(net2768),
    .Y(_06435_));
 NOR2x1_ASAP7_75t_R _12557_ (.A(net2798),
    .B(net2797),
    .Y(_06436_));
 NOR2x1_ASAP7_75t_R _12558_ (.A(net4293),
    .B(_06436_),
    .Y(_06437_));
 OAI21x1_ASAP7_75t_R _12559_ (.A1(_06434_),
    .A2(net2769),
    .B(net2782),
    .Y(_06438_));
 NAND2x1_ASAP7_75t_R _12560_ (.A(_06437_),
    .B(_06438_),
    .Y(_06439_));
 INVx1_ASAP7_75t_R _12561_ (.A(net2770),
    .Y(_06440_));
 NOR2x1_ASAP7_75t_R _12562_ (.A(net2782),
    .B(_06440_),
    .Y(_06441_));
 AOI21x1_ASAP7_75t_R _12563_ (.A1(_06435_),
    .A2(_06439_),
    .B(_06441_),
    .Y(_06442_));
 OAI21x1_ASAP7_75t_R _12564_ (.A1(_06426_),
    .A2(_06425_),
    .B(_06442_),
    .Y(_06443_));
 NOR2x1_ASAP7_75t_R _12565_ (.A(_05438_),
    .B(net4400),
    .Y(_06444_));
 XOR2x2_ASAP7_75t_R _12566_ (.A(_06444_),
    .B(net4721),
    .Y(_06445_));
 AND3x1_ASAP7_75t_R _12567_ (.A(_06445_),
    .B(net4871),
    .C(_05481_),
    .Y(_06446_));
 INVx1_ASAP7_75t_R _12568_ (.A(_06446_),
    .Y(_06447_));
 NOR2x1p5_ASAP7_75t_R _12569_ (.A(net4293),
    .B(_06423_),
    .Y(_06448_));
 INVx1_ASAP7_75t_R _12570_ (.A(net4293),
    .Y(_06449_));
 INVx2_ASAP7_75t_R _12571_ (.A(_06423_),
    .Y(_06450_));
 NOR2x2_ASAP7_75t_R _12572_ (.A(_06450_),
    .B(_06449_),
    .Y(_06451_));
 INVx1_ASAP7_75t_R _12573_ (.A(net2781),
    .Y(_06452_));
 OAI21x1_ASAP7_75t_R _12574_ (.A1(_06448_),
    .A2(_06451_),
    .B(_06452_),
    .Y(_06453_));
 NOR3x1_ASAP7_75t_R _12575_ (.A(_06443_),
    .B(_06447_),
    .C(_06453_),
    .Y(_06454_));
 NAND2x1_ASAP7_75t_R _12576_ (.A(_06423_),
    .B(_06413_),
    .Y(_06455_));
 XOR2x2_ASAP7_75t_R _12577_ (.A(net2783),
    .B(_06455_),
    .Y(_06456_));
 AO21x2_ASAP7_75t_R _12578_ (.A1(_06456_),
    .A2(_06454_),
    .B(net4400),
    .Y(_06457_));
 BUFx3_ASAP7_75t_R place2937 (.A(net5606),
    .Y(net2937));
 BUFx3_ASAP7_75t_R place2936 (.A(_06347_),
    .Y(net2936));
 AO21x1_ASAP7_75t_R _12581_ (.A1(net5114),
    .A2(net5200),
    .B(_06525_),
    .Y(_06460_));
 AOI21x1_ASAP7_75t_R _12582_ (.A1(net5026),
    .A2(net2716),
    .B(_06460_),
    .Y(_00841_));
 AO21x1_ASAP7_75t_R _12583_ (.A1(net2771),
    .A2(_06450_),
    .B(_06425_),
    .Y(_06461_));
 AO21x1_ASAP7_75t_R _12584_ (.A1(_06456_),
    .A2(_06461_),
    .B(net4400),
    .Y(_06462_));
 OA211x2_ASAP7_75t_R _12585_ (.A1(net4871),
    .A2(net4400),
    .B(net4752),
    .C(net5021),
    .Y(_06463_));
 OA21x2_ASAP7_75t_R _12586_ (.A1(net4456),
    .A2(net4664),
    .B(_06463_),
    .Y(_06464_));
 AND2x2_ASAP7_75t_R _12587_ (.A(_06464_),
    .B(_06445_),
    .Y(_06465_));
 OAI21x1_ASAP7_75t_R _12588_ (.A1(_06451_),
    .A2(net2748),
    .B(_06465_),
    .Y(_06466_));
 AO21x1_ASAP7_75t_R _12589_ (.A1(_06423_),
    .A2(_06449_),
    .B(_06452_),
    .Y(_06467_));
 NAND3x1_ASAP7_75t_R _12590_ (.A(_06467_),
    .B(_06442_),
    .C(net2750),
    .Y(_06468_));
 OAI21x1_ASAP7_75t_R _12591_ (.A1(_06468_),
    .A2(_06466_),
    .B(net4456),
    .Y(_06469_));
 AND2x4_ASAP7_75t_R _12592_ (.A(_06469_),
    .B(_06462_),
    .Y(_06470_));
 BUFx3_ASAP7_75t_R place2934 (.A(_04002_),
    .Y(net2934));
 BUFx3_ASAP7_75t_R place2933 (.A(_04002_),
    .Y(net2933));
 AO21x1_ASAP7_75t_R _12595_ (.A1(net5113),
    .A2(net5200),
    .B(_06525_),
    .Y(_06473_));
 AOI21x1_ASAP7_75t_R _12596_ (.A1(net5026),
    .A2(net2715),
    .B(_06473_),
    .Y(_00842_));
 AO21x1_ASAP7_75t_R _12597_ (.A1(net5112),
    .A2(net5200),
    .B(_06525_),
    .Y(_06474_));
 AOI21x1_ASAP7_75t_R _12598_ (.A1(net5026),
    .A2(net2716),
    .B(_06474_),
    .Y(_00843_));
 AO21x1_ASAP7_75t_R _12599_ (.A1(net5111),
    .A2(net5200),
    .B(_06525_),
    .Y(_06475_));
 AOI21x1_ASAP7_75t_R _12600_ (.A1(net5026),
    .A2(net2715),
    .B(_06475_),
    .Y(_00844_));
 BUFx6f_ASAP7_75t_R place2932 (.A(_05187_),
    .Y(net2932));
 AO21x1_ASAP7_75t_R _12602_ (.A1(net5110),
    .A2(net5200),
    .B(_06525_),
    .Y(_06477_));
 AOI21x1_ASAP7_75t_R _12603_ (.A1(net5024),
    .A2(net2716),
    .B(_06477_),
    .Y(_00845_));
 AO21x1_ASAP7_75t_R _12604_ (.A1(net5109),
    .A2(net5200),
    .B(_06525_),
    .Y(_06478_));
 AOI21x1_ASAP7_75t_R _12605_ (.A1(net5026),
    .A2(net2715),
    .B(_06478_),
    .Y(_00846_));
 AO21x1_ASAP7_75t_R _12606_ (.A1(net5108),
    .A2(net5200),
    .B(_06525_),
    .Y(_06479_));
 AOI21x1_ASAP7_75t_R _12607_ (.A1(net2717),
    .A2(net5026),
    .B(_06479_),
    .Y(_00847_));
 AO21x1_ASAP7_75t_R _12608_ (.A1(net5107),
    .A2(net5200),
    .B(_06525_),
    .Y(_06480_));
 AOI21x1_ASAP7_75t_R _12609_ (.A1(net5026),
    .A2(net2715),
    .B(_06480_),
    .Y(_00848_));
 AO21x1_ASAP7_75t_R _12610_ (.A1(net5106),
    .A2(net5200),
    .B(_06525_),
    .Y(_06481_));
 AOI21x1_ASAP7_75t_R _12611_ (.A1(net5026),
    .A2(net2716),
    .B(_06481_),
    .Y(_00849_));
 AO21x1_ASAP7_75t_R _12612_ (.A1(net5105),
    .A2(net5200),
    .B(_06525_),
    .Y(_06482_));
 AOI21x1_ASAP7_75t_R _12613_ (.A1(net2714),
    .A2(net5025),
    .B(_06482_),
    .Y(_00850_));
 BUFx3_ASAP7_75t_R place2930 (.A(_05203_),
    .Y(net2930));
 AO21x1_ASAP7_75t_R _12615_ (.A1(net5200),
    .A2(net5104),
    .B(_06525_),
    .Y(_06484_));
 AOI21x1_ASAP7_75t_R _12616_ (.A1(net5027),
    .A2(net4752),
    .B(_06484_),
    .Y(_00851_));
 BUFx3_ASAP7_75t_R place2929 (.A(_05240_),
    .Y(net2929));
 AO21x1_ASAP7_75t_R _12618_ (.A1(net5103),
    .A2(net5200),
    .B(_06525_),
    .Y(_06486_));
 AOI21x1_ASAP7_75t_R _12619_ (.A1(net2717),
    .A2(net5025),
    .B(_06486_),
    .Y(_00852_));
 AO21x1_ASAP7_75t_R _12620_ (.A1(net5102),
    .A2(net5200),
    .B(_06525_),
    .Y(_06487_));
 AOI21x1_ASAP7_75t_R _12621_ (.A1(net5025),
    .A2(net2714),
    .B(_06487_),
    .Y(_00853_));
 AO21x1_ASAP7_75t_R _12622_ (.A1(net5101),
    .A2(net5200),
    .B(_06525_),
    .Y(_06488_));
 AOI21x1_ASAP7_75t_R _12623_ (.A1(net2717),
    .A2(net5025),
    .B(_06488_),
    .Y(_00854_));
 AO21x1_ASAP7_75t_R _12624_ (.A1(net5100),
    .A2(net5200),
    .B(_06525_),
    .Y(_06489_));
 AOI21x1_ASAP7_75t_R _12625_ (.A1(net5025),
    .A2(net2714),
    .B(_06489_),
    .Y(_00855_));
 BUFx3_ASAP7_75t_R place2931 (.A(net2930),
    .Y(net2931));
 AO21x1_ASAP7_75t_R _12627_ (.A1(net5099),
    .A2(net5200),
    .B(_06525_),
    .Y(_06491_));
 AOI21x1_ASAP7_75t_R _12628_ (.A1(net2717),
    .A2(net5025),
    .B(_06491_),
    .Y(_00856_));
 AO21x1_ASAP7_75t_R _12629_ (.A1(net5098),
    .A2(net5200),
    .B(_06525_),
    .Y(_06492_));
 AOI21x1_ASAP7_75t_R _12630_ (.A1(net5025),
    .A2(net2714),
    .B(_06492_),
    .Y(_00857_));
 AO21x1_ASAP7_75t_R _12631_ (.A1(net5096),
    .A2(net5200),
    .B(_06525_),
    .Y(_06493_));
 AOI21x1_ASAP7_75t_R _12632_ (.A1(net2717),
    .A2(net5025),
    .B(_06493_),
    .Y(_00858_));
 AO21x1_ASAP7_75t_R _12633_ (.A1(net5095),
    .A2(net5200),
    .B(_06525_),
    .Y(_06494_));
 AOI21x1_ASAP7_75t_R _12634_ (.A1(net2714),
    .A2(net5025),
    .B(_06494_),
    .Y(_00859_));
 AO21x1_ASAP7_75t_R _12635_ (.A1(_00050_),
    .A2(net5200),
    .B(_06525_),
    .Y(_06495_));
 AOI21x1_ASAP7_75t_R _12636_ (.A1(net2717),
    .A2(net5025),
    .B(_06495_),
    .Y(_00860_));
 AO21x1_ASAP7_75t_R _12637_ (.A1(net5094),
    .A2(net5200),
    .B(_06525_),
    .Y(_06496_));
 AOI21x1_ASAP7_75t_R _12638_ (.A1(net2714),
    .A2(net5025),
    .B(_06496_),
    .Y(_00861_));
 OA21x2_ASAP7_75t_R _12639_ (.A1(net4871),
    .A2(net5024),
    .B(net5363),
    .Y(_06497_));
 OA21x2_ASAP7_75t_R _12640_ (.A1(net5200),
    .A2(net4720),
    .B(_06497_),
    .Y(_00862_));
 AO21x1_ASAP7_75t_R _12641_ (.A1(net5091),
    .A2(net5200),
    .B(_06525_),
    .Y(_06498_));
 AOI21x1_ASAP7_75t_R _12642_ (.A1(net2717),
    .A2(net5025),
    .B(_06498_),
    .Y(_00863_));
 AO21x1_ASAP7_75t_R _12643_ (.A1(net5090),
    .A2(net5200),
    .B(_06525_),
    .Y(_06499_));
 AOI21x1_ASAP7_75t_R _12644_ (.A1(net5026),
    .A2(net2714),
    .B(_06499_),
    .Y(_00864_));
 NOR2x1p5_ASAP7_75t_R _12645_ (.A(net4400),
    .B(net4291),
    .Y(_06500_));
 XOR2x2_ASAP7_75t_R _12646_ (.A(net4292),
    .B(_06500_),
    .Y(_06501_));
 AO21x1_ASAP7_75t_R _12647_ (.A1(net5200),
    .A2(net5089),
    .B(_06525_),
    .Y(_06502_));
 AOI21x1_ASAP7_75t_R _12648_ (.A1(net5027),
    .A2(_06501_),
    .B(_06502_),
    .Y(_00865_));
 NOR2x2_ASAP7_75t_R _12649_ (.A(net2740),
    .B(net5957),
    .Y(_06503_));
 NAND2x1_ASAP7_75t_R _12650_ (.A(net4456),
    .B(_06447_),
    .Y(_06504_));
 XOR2x2_ASAP7_75t_R _12651_ (.A(_06503_),
    .B(_06504_),
    .Y(_06505_));
 AO21x1_ASAP7_75t_R _12652_ (.A1(net5088),
    .A2(net5200),
    .B(_06525_),
    .Y(_06506_));
 AOI21x1_ASAP7_75t_R _12653_ (.A1(net5027),
    .A2(_06505_),
    .B(_06506_),
    .Y(_00866_));
 NAND2x1_ASAP7_75t_R _12654_ (.A(net4456),
    .B(net5662),
    .Y(_06507_));
 AND2x2_ASAP7_75t_R _12655_ (.A(_06467_),
    .B(net2750),
    .Y(_06508_));
 XOR2x2_ASAP7_75t_R _12656_ (.A(_06507_),
    .B(_06508_),
    .Y(_06509_));
 OA21x2_ASAP7_75t_R _12657_ (.A1(net5012),
    .A2(net5024),
    .B(net5363),
    .Y(_06510_));
 OA21x2_ASAP7_75t_R _12658_ (.A1(_06509_),
    .A2(net5200),
    .B(_06510_),
    .Y(_00867_));
 OA21x2_ASAP7_75t_R _12659_ (.A1(net2733),
    .A2(_06447_),
    .B(net4456),
    .Y(_06511_));
 XOR2x2_ASAP7_75t_R _12660_ (.A(_06511_),
    .B(net2741),
    .Y(_06512_));
 AO21x1_ASAP7_75t_R _12661_ (.A1(net5086),
    .A2(net5200),
    .B(_06525_),
    .Y(_06513_));
 AOI21x1_ASAP7_75t_R _12662_ (.A1(net5027),
    .A2(_06512_),
    .B(_06513_),
    .Y(_00868_));
 INVx1_ASAP7_75t_R _12663_ (.A(net2727),
    .Y(_06514_));
 AOI21x1_ASAP7_75t_R _12664_ (.A1(_06514_),
    .A2(net5661),
    .B(net5200),
    .Y(_06515_));
 OR2x2_ASAP7_75t_R _12665_ (.A(_06514_),
    .B(net5661),
    .Y(_06516_));
 AO21x1_ASAP7_75t_R _12666_ (.A1(net5085),
    .A2(net5200),
    .B(_06525_),
    .Y(_06517_));
 AOI21x1_ASAP7_75t_R _12667_ (.A1(_06515_),
    .A2(_06516_),
    .B(_06517_),
    .Y(_00869_));
 OAI21x1_ASAP7_75t_R _12668_ (.A1(net2733),
    .A2(net5653),
    .B(net4456),
    .Y(_06518_));
 INVx1_ASAP7_75t_R _12669_ (.A(net2739),
    .Y(_06519_));
 NAND3x1_ASAP7_75t_R _12670_ (.A(_06518_),
    .B(_06519_),
    .C(net4105),
    .Y(_06520_));
 NAND2x1_ASAP7_75t_R _12671_ (.A(_06504_),
    .B(_06518_),
    .Y(_06521_));
 AOI21x1_ASAP7_75t_R _12672_ (.A1(net2739),
    .A2(_06521_),
    .B(net5200),
    .Y(_06522_));
 AO21x1_ASAP7_75t_R _12673_ (.A1(net5084),
    .A2(net5200),
    .B(_06525_),
    .Y(_06523_));
 AOI21x1_ASAP7_75t_R _12674_ (.A1(_06522_),
    .A2(_06520_),
    .B(_06523_),
    .Y(_00870_));
 AO21x1_ASAP7_75t_R _12675_ (.A1(net5083),
    .A2(net5200),
    .B(_06525_),
    .Y(_06524_));
 AOI21x1_ASAP7_75t_R _12676_ (.A1(net5026),
    .A2(net2715),
    .B(_06524_),
    .Y(_00871_));
 INVx1_ASAP7_75t_R _12677_ (.A(_00368_),
    .Y(_00369_));
 FAx1_ASAP7_75t_R _12678_ (.SN(_00340_),
    .A(net5071),
    .B(net4927),
    .CI(_00338_),
    .CON(_00339_));
 HAxp5_ASAP7_75t_R _12679_ (.A(\u_fft.sched[54] ),
    .B(_00341_),
    .CON(_00342_),
    .SN(_00343_));
 HAxp5_ASAP7_75t_R _12680_ (.A(_00344_),
    .B(\u_fft.sched[53] ),
    .CON(_00345_),
    .SN(_00346_));
 HAxp5_ASAP7_75t_R _12681_ (.A(\u_fft.sched[52] ),
    .B(_00347_),
    .CON(_00348_),
    .SN(_00349_));
 HAxp5_ASAP7_75t_R _12682_ (.A(\u_fft.sched[51] ),
    .B(_00350_),
    .CON(_00351_),
    .SN(_00352_));
 HAxp5_ASAP7_75t_R _12683_ (.A(_00353_),
    .B(\u_fft.sched[50] ),
    .CON(_00354_),
    .SN(_00355_));
 HAxp5_ASAP7_75t_R _12684_ (.A(\u_fft.sched[49] ),
    .B(_00356_),
    .CON(_00357_),
    .SN(_00358_));
 HAxp5_ASAP7_75t_R _12685_ (.A(\u_fft.sched[48] ),
    .B(_00359_),
    .CON(_00360_),
    .SN(_00361_));
 HAxp5_ASAP7_75t_R _12686_ (.A(\u_fft.sched[47] ),
    .B(_00362_),
    .CON(_00363_),
    .SN(_00364_));
 HAxp5_ASAP7_75t_R _12687_ (.A(_00366_),
    .B(_00365_),
    .CON(_00367_),
    .SN(_00368_));
 HAxp5_ASAP7_75t_R _12688_ (.A(\u_fft.sched[46] ),
    .B(_00369_),
    .CON(_00370_),
    .SN(_00371_));
 HAxp5_ASAP7_75t_R _12689_ (.A(\u_fft.sched[64] ),
    .B(_00372_),
    .CON(_00373_),
    .SN(_00374_));
 HAxp5_ASAP7_75t_R _12690_ (.A(\u_fft.sched[63] ),
    .B(_00375_),
    .CON(_00376_),
    .SN(_00377_));
 HAxp5_ASAP7_75t_R _12691_ (.A(\u_fft.sched[62] ),
    .B(_00378_),
    .CON(_00379_),
    .SN(_00380_));
 HAxp5_ASAP7_75t_R _12692_ (.A(\u_fft.sched[61] ),
    .B(_00381_),
    .CON(_00382_),
    .SN(_00383_));
 HAxp5_ASAP7_75t_R _12693_ (.A(\u_fft.sched[60] ),
    .B(_00384_),
    .CON(_00385_),
    .SN(_00386_));
 HAxp5_ASAP7_75t_R _12694_ (.A(\u_fft.sched[59] ),
    .B(_00387_),
    .CON(_00388_),
    .SN(_00389_));
 HAxp5_ASAP7_75t_R _12695_ (.A(\u_fft.sched[58] ),
    .B(_00390_),
    .CON(_00391_),
    .SN(_00392_));
 HAxp5_ASAP7_75t_R _12696_ (.A(\u_fft.sched[57] ),
    .B(_00393_),
    .CON(_00394_),
    .SN(_00395_));
 HAxp5_ASAP7_75t_R _12697_ (.A(net5273),
    .B(_00397_),
    .CON(_00398_),
    .SN(_06529_));
 HAxp5_ASAP7_75t_R _12698_ (.A(\u_fft.sched[56] ),
    .B(_06529_),
    .CON(_00399_),
    .SN(_00400_));
 HAxp5_ASAP7_75t_R _12699_ (.A(\u_window_buffer.read_ptr[30] ),
    .B(\u_window_buffer.internal_read_ptr[30] ),
    .CON(_00401_),
    .SN(_00402_));
 HAxp5_ASAP7_75t_R _12700_ (.A(\u_window_buffer.read_ptr[29] ),
    .B(\u_window_buffer.internal_read_ptr[29] ),
    .CON(_00403_),
    .SN(_00404_));
 HAxp5_ASAP7_75t_R _12701_ (.A(\u_window_buffer.read_ptr[28] ),
    .B(\u_window_buffer.internal_read_ptr[28] ),
    .CON(_00405_),
    .SN(_00406_));
 HAxp5_ASAP7_75t_R _12702_ (.A(\u_window_buffer.internal_read_ptr[27] ),
    .B(\u_window_buffer.read_ptr[27] ),
    .CON(_00407_),
    .SN(_00408_));
 HAxp5_ASAP7_75t_R _12703_ (.A(\u_window_buffer.read_ptr[26] ),
    .B(\u_window_buffer.internal_read_ptr[26] ),
    .CON(_00409_),
    .SN(_00410_));
 HAxp5_ASAP7_75t_R _12704_ (.A(\u_window_buffer.read_ptr[25] ),
    .B(\u_window_buffer.internal_read_ptr[25] ),
    .CON(_00411_),
    .SN(_00412_));
 HAxp5_ASAP7_75t_R _12705_ (.A(\u_window_buffer.internal_read_ptr[24] ),
    .B(\u_window_buffer.read_ptr[24] ),
    .CON(_00413_),
    .SN(_00414_));
 HAxp5_ASAP7_75t_R _12706_ (.A(\u_window_buffer.internal_read_ptr[23] ),
    .B(\u_window_buffer.read_ptr[23] ),
    .CON(_00415_),
    .SN(_00416_));
 HAxp5_ASAP7_75t_R _12707_ (.A(\u_window_buffer.read_ptr[22] ),
    .B(\u_window_buffer.internal_read_ptr[22] ),
    .CON(_00417_),
    .SN(_00418_));
 HAxp5_ASAP7_75t_R _12708_ (.A(\u_window_buffer.read_ptr[21] ),
    .B(\u_window_buffer.internal_read_ptr[21] ),
    .CON(_00419_),
    .SN(_00420_));
 HAxp5_ASAP7_75t_R _12709_ (.A(\u_window_buffer.read_ptr[20] ),
    .B(\u_window_buffer.internal_read_ptr[20] ),
    .CON(_00421_),
    .SN(_00422_));
 HAxp5_ASAP7_75t_R _12710_ (.A(\u_window_buffer.read_ptr[19] ),
    .B(\u_window_buffer.internal_read_ptr[19] ),
    .CON(_00423_),
    .SN(_00424_));
 HAxp5_ASAP7_75t_R _12711_ (.A(\u_window_buffer.internal_read_ptr[18] ),
    .B(\u_window_buffer.read_ptr[18] ),
    .CON(_00425_),
    .SN(_00426_));
 HAxp5_ASAP7_75t_R _12712_ (.A(\u_window_buffer.read_ptr[17] ),
    .B(\u_window_buffer.internal_read_ptr[17] ),
    .CON(_00427_),
    .SN(_00428_));
 HAxp5_ASAP7_75t_R _12713_ (.A(\u_window_buffer.internal_read_ptr[16] ),
    .B(\u_window_buffer.read_ptr[16] ),
    .CON(_00429_),
    .SN(_00430_));
 HAxp5_ASAP7_75t_R _12714_ (.A(\u_window_buffer.read_ptr[15] ),
    .B(\u_window_buffer.internal_read_ptr[15] ),
    .CON(_00431_),
    .SN(_00432_));
 HAxp5_ASAP7_75t_R _12715_ (.A(\u_window_buffer.internal_read_ptr[14] ),
    .B(\u_window_buffer.read_ptr[14] ),
    .CON(_00433_),
    .SN(_00434_));
 HAxp5_ASAP7_75t_R _12716_ (.A(\u_window_buffer.internal_read_ptr[13] ),
    .B(\u_window_buffer.read_ptr[13] ),
    .CON(_00435_),
    .SN(_00436_));
 HAxp5_ASAP7_75t_R _12717_ (.A(\u_window_buffer.read_ptr[12] ),
    .B(\u_window_buffer.internal_read_ptr[12] ),
    .CON(_00437_),
    .SN(_00438_));
 HAxp5_ASAP7_75t_R _12718_ (.A(\u_window_buffer.internal_read_ptr[11] ),
    .B(\u_window_buffer.read_ptr[11] ),
    .CON(_00439_),
    .SN(_00440_));
 HAxp5_ASAP7_75t_R _12719_ (.A(\u_window_buffer.internal_read_ptr[10] ),
    .B(\u_window_buffer.read_ptr[10] ),
    .CON(_00441_),
    .SN(_00442_));
 HAxp5_ASAP7_75t_R _12720_ (.A(\u_window_buffer.read_ptr[9] ),
    .B(\u_window_buffer.internal_read_ptr[9] ),
    .CON(_00443_),
    .SN(_00444_));
 HAxp5_ASAP7_75t_R _12721_ (.A(\u_window_buffer.read_ptr[8] ),
    .B(\u_window_buffer.internal_read_ptr[8] ),
    .CON(_00445_),
    .SN(_00446_));
 HAxp5_ASAP7_75t_R _12722_ (.A(\u_window_buffer.internal_read_ptr[7] ),
    .B(\u_window_buffer.read_ptr[7] ),
    .CON(_00447_),
    .SN(_00448_));
 HAxp5_ASAP7_75t_R _12723_ (.A(\u_window_buffer.internal_read_ptr[6] ),
    .B(\u_window_buffer.read_ptr[6] ),
    .CON(_00449_),
    .SN(_00450_));
 HAxp5_ASAP7_75t_R _12724_ (.A(\u_window_buffer.read_ptr[5] ),
    .B(\u_window_buffer.internal_read_ptr[5] ),
    .CON(_00451_),
    .SN(_00452_));
 HAxp5_ASAP7_75t_R _12725_ (.A(\u_window_buffer.read_ptr[4] ),
    .B(\u_window_buffer.internal_read_ptr[4] ),
    .CON(_00453_),
    .SN(_00454_));
 HAxp5_ASAP7_75t_R _12726_ (.A(\u_window_buffer.read_ptr[3] ),
    .B(\u_window_buffer.internal_read_ptr[3] ),
    .CON(_00455_),
    .SN(_00456_));
 HAxp5_ASAP7_75t_R _12727_ (.A(\u_window_buffer.read_ptr[2] ),
    .B(\u_window_buffer.internal_read_ptr[2] ),
    .CON(_00457_),
    .SN(_00458_));
 HAxp5_ASAP7_75t_R _12728_ (.A(net4935),
    .B(\u_window_buffer.internal_read_ptr[1] ),
    .CON(_00459_),
    .SN(_00462_));
 HAxp5_ASAP7_75t_R _12729_ (.A(net4935),
    .B(\u_window_buffer.internal_read_ptr[1] ),
    .CON(_00460_),
    .SN(_06530_));
 HAxp5_ASAP7_75t_R _12730_ (.A(net5143),
    .B(net4760),
    .CON(_00463_),
    .SN(_00464_));
 HAxp5_ASAP7_75t_R _12731_ (.A(net5143),
    .B(_00465_),
    .CON(_00466_),
    .SN(_00467_));
 HAxp5_ASAP7_75t_R _12732_ (.A(\tx_fifo.write_ptr[1] ),
    .B(\tx_fifo.write_ptr[0] ),
    .CON(_00468_),
    .SN(_00469_));
 HAxp5_ASAP7_75t_R _12733_ (.A(_00470_),
    .B(_00471_),
    .CON(_00472_),
    .SN(_00473_));
 HAxp5_ASAP7_75t_R _12734_ (.A(\u_dct.k_ptr[0] ),
    .B(\u_dct.k_ptr[1] ),
    .CON(_00474_),
    .SN(_06531_));
 HAxp5_ASAP7_75t_R _12735_ (.A(net5337),
    .B(net5336),
    .CON(_00477_),
    .SN(_00478_));
 HAxp5_ASAP7_75t_R _12736_ (.A(\u_dct.n_ptr[0] ),
    .B(\u_dct.n_ptr[1] ),
    .CON(_00479_),
    .SN(_06532_));
 HAxp5_ASAP7_75t_R _12737_ (.A(net5264),
    .B(net5263),
    .CON(_00482_),
    .SN(_00483_));
 HAxp5_ASAP7_75t_R _12738_ (.A(net5264),
    .B(net5067),
    .CON(_00484_),
    .SN(_06533_));
 HAxp5_ASAP7_75t_R _12739_ (.A(net5066),
    .B(net5263),
    .CON(_00485_),
    .SN(_06534_));
 HAxp5_ASAP7_75t_R _12740_ (.A(\u_fft.sched[40] ),
    .B(\u_fft.sched[41] ),
    .CON(_00486_),
    .SN(_06535_));
 HAxp5_ASAP7_75t_R _12741_ (.A(net5262),
    .B(_00487_),
    .CON(_00489_),
    .SN(_00490_));
 HAxp5_ASAP7_75t_R _12742_ (.A(net5068),
    .B(net4745),
    .CON(_00491_),
    .SN(_06536_));
 HAxp5_ASAP7_75t_R _12743_ (.A(\u_fft.sched[45] ),
    .B(net4999),
    .CON(_00492_),
    .SN(_00493_));
 HAxp5_ASAP7_75t_R _12744_ (.A(net5070),
    .B(_00494_),
    .CON(_00495_),
    .SN(_00496_));
 HAxp5_ASAP7_75t_R _12745_ (.A(net5070),
    .B(\u_fft.sched[55] ),
    .CON(_00497_),
    .SN(_06537_));
 HAxp5_ASAP7_75t_R _12746_ (.A(net5071),
    .B(net4927),
    .CON(_00498_),
    .SN(_00499_));
 HAxp5_ASAP7_75t_R _12747_ (.A(net5072),
    .B(\u_fft.sched[57] ),
    .CON(_00500_),
    .SN(_00501_));
 HAxp5_ASAP7_75t_R _12748_ (.A(net5073),
    .B(net4928),
    .CON(_00502_),
    .SN(_00503_));
 HAxp5_ASAP7_75t_R _12749_ (.A(net5074),
    .B(net4929),
    .CON(_00504_),
    .SN(_00505_));
 HAxp5_ASAP7_75t_R _12750_ (.A(net5075),
    .B(net4930),
    .CON(_00506_),
    .SN(_00507_));
 HAxp5_ASAP7_75t_R _12751_ (.A(net5076),
    .B(net4931),
    .CON(_00508_),
    .SN(_00509_));
 HAxp5_ASAP7_75t_R _12752_ (.A(net5077),
    .B(\u_fft.sched[62] ),
    .CON(_00510_),
    .SN(_00511_));
 HAxp5_ASAP7_75t_R _12753_ (.A(net5078),
    .B(net4932),
    .CON(_00512_),
    .SN(_00513_));
 HAxp5_ASAP7_75t_R _12754_ (.A(\u_fft.power_ptr[0] ),
    .B(\u_fft.power_ptr[1] ),
    .CON(_00514_),
    .SN(_00515_));
 HAxp5_ASAP7_75t_R _12755_ (.A(\u_hamming_window.frame_ptr[0] ),
    .B(\u_hamming_window.frame_ptr[1] ),
    .CON(_00516_),
    .SN(_00517_));
 HAxp5_ASAP7_75t_R _12756_ (.A(_00519_),
    .B(_00518_),
    .CON(_00520_),
    .SN(_00521_));
 HAxp5_ASAP7_75t_R _12757_ (.A(\mel_ptr[0] ),
    .B(\mel_ptr[1] ),
    .CON(_00522_),
    .SN(_06538_));
 HAxp5_ASAP7_75t_R _12758_ (.A(net5189),
    .B(net5179),
    .CON(_00525_),
    .SN(_00526_));
 HAxp5_ASAP7_75t_R _12759_ (.A(net5189),
    .B(net5179),
    .CON(_00527_),
    .SN(_06539_));
 HAxp5_ASAP7_75t_R _12760_ (.A(net5189),
    .B(_00528_),
    .CON(_00529_),
    .SN(_00530_));
 HAxp5_ASAP7_75t_R _12761_ (.A(net5709),
    .B(net4964),
    .CON(_00531_),
    .SN(_00532_));
 HAxp5_ASAP7_75t_R _12762_ (.A(net4965),
    .B(net4964),
    .CON(_00533_),
    .SN(_06540_));
 HAxp5_ASAP7_75t_R _12763_ (.A(net5163),
    .B(net5171),
    .CON(_00536_),
    .SN(_00537_));
 HAxp5_ASAP7_75t_R _12764_ (.A(\u_window_buffer.move_counter[0] ),
    .B(net5163),
    .CON(_00538_),
    .SN(_06541_));
 HAxp5_ASAP7_75t_R _12765_ (.A(\u_window_buffer.read_ptr[0] ),
    .B(\u_window_buffer.read_ptr[1] ),
    .CON(_00539_),
    .SN(_00540_));
 HAxp5_ASAP7_75t_R _12766_ (.A(\u_window_buffer.write_ptr[0] ),
    .B(\u_window_buffer.write_ptr[1] ),
    .CON(_00541_),
    .SN(_00542_));
 HAxp5_ASAP7_75t_R _12767_ (.A(net5357),
    .B(net5356),
    .CON(_00545_),
    .SN(_00546_));
 HAxp5_ASAP7_75t_R _12768_ (.A(\tx_fifo.read_ptr[0] ),
    .B(\tx_fifo.read_ptr[1] ),
    .CON(_00547_),
    .SN(_06542_));
 HAxp5_ASAP7_75t_R _12769_ (.A(net5241),
    .B(net5249),
    .CON(_00550_),
    .SN(_00551_));
 HAxp5_ASAP7_75t_R _12770_ (.A(\u_hamming_window.calc_pointer[0] ),
    .B(\u_hamming_window.calc_pointer[1] ),
    .CON(_00552_),
    .SN(_06543_));
 HAxp5_ASAP7_75t_R _12771_ (.A(_00553_),
    .B(\u_mel.k_next[0] ),
    .CON(_00554_),
    .SN(_00555_));
 HAxp5_ASAP7_75t_R _12772_ (.A(\u_mel.k[0] ),
    .B(\u_mel.k[1] ),
    .CON(_00556_),
    .SN(_06544_));
 DFFHQNx1_ASAP7_75t_R _12773_ (.CLK(clknet_leaf_20_clk),
    .D(_00021_),
    .QN(_00054_));
 DFFHQNx1_ASAP7_75t_R _12774_ (.CLK(clknet_leaf_20_clk),
    .D(_00022_),
    .QN(_00056_));
 BUFx3_ASAP7_75t_R place2928 (.A(_05274_),
    .Y(net2928));
 BUFx3_ASAP7_75t_R place2927 (.A(_06318_),
    .Y(net2927));
 BUFx3_ASAP7_75t_R place2926 (.A(_02257_),
    .Y(net2926));
 BUFx3_ASAP7_75t_R place2924 (.A(net5447),
    .Y(net2924));
 BUFx3_ASAP7_75t_R place2923 (.A(_02301_),
    .Y(net2923));
 BUFx3_ASAP7_75t_R place2921 (.A(_04011_),
    .Y(net2921));
 BUFx3_ASAP7_75t_R place2920 (.A(_04012_),
    .Y(net2920));
 BUFx3_ASAP7_75t_R place2918 (.A(net5620),
    .Y(net2918));
 BUFx3_ASAP7_75t_R place2919 (.A(_05219_),
    .Y(net2919));
 BUFx3_ASAP7_75t_R place2917 (.A(_06354_),
    .Y(net2917));
 BUFx3_ASAP7_75t_R place2916 (.A(_02286_),
    .Y(net2916));
 BUFx3_ASAP7_75t_R place2915 (.A(net5391),
    .Y(net2915));
 BUFx3_ASAP7_75t_R place2914 (.A(_02297_),
    .Y(net2914));
 BUFx3_ASAP7_75t_R place2912 (.A(_02306_),
    .Y(net2912));
 BUFx3_ASAP7_75t_R place2911 (.A(_02315_),
    .Y(net2911));
 BUFx3_ASAP7_75t_R place2910 (.A(_02316_),
    .Y(net2910));
 BUFx3_ASAP7_75t_R place2908 (.A(_03995_),
    .Y(net2908));
 BUFx3_ASAP7_75t_R place2907 (.A(_04005_),
    .Y(net2907));
 BUFx3_ASAP7_75t_R place2906 (.A(_04013_),
    .Y(net2906));
 BUFx3_ASAP7_75t_R place2905 (.A(_04017_),
    .Y(net2905));
 BUFx3_ASAP7_75t_R place2904 (.A(_04024_),
    .Y(net2904));
 BUFx3_ASAP7_75t_R place2903 (.A(_04030_),
    .Y(net2903));
 BUFx3_ASAP7_75t_R place2902 (.A(_05242_),
    .Y(net2902));
 BUFx3_ASAP7_75t_R place2901 (.A(_05243_),
    .Y(net2901));
 BUFx3_ASAP7_75t_R place2909 (.A(_03990_),
    .Y(net2909));
 BUFx6f_ASAP7_75t_R place2900 (.A(_05247_),
    .Y(net2900));
 BUFx3_ASAP7_75t_R place2898 (.A(_06338_),
    .Y(net2898));
 BUFx3_ASAP7_75t_R place2897 (.A(_06340_),
    .Y(net2897));
 BUFx3_ASAP7_75t_R place2896 (.A(_06355_),
    .Y(net2896));
 BUFx3_ASAP7_75t_R place2895 (.A(_06379_),
    .Y(net2895));
 BUFx3_ASAP7_75t_R place2894 (.A(_06384_),
    .Y(net2894));
 BUFx3_ASAP7_75t_R place2893 (.A(_02280_),
    .Y(net2893));
 BUFx3_ASAP7_75t_R place2892 (.A(_02280_),
    .Y(net2892));
 BUFx3_ASAP7_75t_R place2888 (.A(_02317_),
    .Y(net2888));
 BUFx3_ASAP7_75t_R place2887 (.A(net5537),
    .Y(net2887));
 BUFx3_ASAP7_75t_R place2886 (.A(_03996_),
    .Y(net2886));
 BUFx3_ASAP7_75t_R place2885 (.A(_04014_),
    .Y(net2885));
 BUFx3_ASAP7_75t_R place2884 (.A(net5684),
    .Y(net2884));
 BUFx3_ASAP7_75t_R place2883 (.A(_05244_),
    .Y(net2883));
 BUFx3_ASAP7_75t_R place2882 (.A(_06334_),
    .Y(net2882));
 BUFx3_ASAP7_75t_R place2880 (.A(_06362_),
    .Y(net2880));
 BUFx3_ASAP7_75t_R place2878 (.A(_06382_),
    .Y(net2878));
 BUFx3_ASAP7_75t_R place2877 (.A(_02308_),
    .Y(net2877));
 BUFx3_ASAP7_75t_R place2874 (.A(_04026_),
    .Y(net2874));
 BUFx3_ASAP7_75t_R place2873 (.A(_04035_),
    .Y(net2873));
 BUFx3_ASAP7_75t_R place2872 (.A(_05224_),
    .Y(net2872));
 BUFx3_ASAP7_75t_R place2871 (.A(_05246_),
    .Y(net2871));
 BUFx3_ASAP7_75t_R place2869 (.A(_05263_),
    .Y(net2869));
 BUFx3_ASAP7_75t_R place2870 (.A(_05248_),
    .Y(net2870));
 BUFx6f_ASAP7_75t_R place2867 (.A(_06341_),
    .Y(net2867));
 BUFx3_ASAP7_75t_R place2865 (.A(_06356_),
    .Y(net2865));
 BUFx3_ASAP7_75t_R place2864 (.A(_02289_),
    .Y(net2864));
 BUFx3_ASAP7_75t_R place2866 (.A(_06349_),
    .Y(net2866));
 BUFx3_ASAP7_75t_R place2863 (.A(net5821),
    .Y(net2863));
 BUFx6f_ASAP7_75t_R place2862 (.A(_02332_),
    .Y(net2862));
 BUFx3_ASAP7_75t_R place2861 (.A(_02336_),
    .Y(net2861));
 BUFx3_ASAP7_75t_R place2860 (.A(_02339_),
    .Y(net2860));
 BUFx3_ASAP7_75t_R place2859 (.A(_02352_),
    .Y(net2859));
 BUFx3_ASAP7_75t_R place2868 (.A(net2867),
    .Y(net2868));
 BUFx3_ASAP7_75t_R place2858 (.A(_04036_),
    .Y(net2858));
 BUFx3_ASAP7_75t_R place2857 (.A(_04038_),
    .Y(net2857));
 BUFx3_ASAP7_75t_R place2854 (.A(_05250_),
    .Y(net2854));
 BUFx3_ASAP7_75t_R place2853 (.A(_05259_),
    .Y(net2853));
 BUFx3_ASAP7_75t_R place2852 (.A(_05264_),
    .Y(net2852));
 BUFx3_ASAP7_75t_R place2855 (.A(_05225_),
    .Y(net2855));
 BUFx3_ASAP7_75t_R place2851 (.A(_05273_),
    .Y(net2851));
 BUFx3_ASAP7_75t_R place2856 (.A(_04046_),
    .Y(net2856));
 BUFx3_ASAP7_75t_R place2850 (.A(_05285_),
    .Y(net2850));
 BUFx3_ASAP7_75t_R place2849 (.A(net5618),
    .Y(net2849));
 BUFx3_ASAP7_75t_R place2848 (.A(_06369_),
    .Y(net2848));
 BUFx3_ASAP7_75t_R place2847 (.A(_02300_),
    .Y(net2847));
 BUFx3_ASAP7_75t_R place2846 (.A(_02333_),
    .Y(net2846));
 BUFx3_ASAP7_75t_R place2875 (.A(_04000_),
    .Y(net2875));
 BUFx3_ASAP7_75t_R place2843 (.A(_04019_),
    .Y(net2843));
 BUFx3_ASAP7_75t_R place2842 (.A(_04044_),
    .Y(net2842));
 BUFx3_ASAP7_75t_R place2841 (.A(_04056_),
    .Y(net2841));
 BUFx3_ASAP7_75t_R place2840 (.A(_04060_),
    .Y(net2840));
 BUFx3_ASAP7_75t_R place2838 (.A(_05254_),
    .Y(net2838));
 BUFx3_ASAP7_75t_R place2836 (.A(net5614),
    .Y(net2836));
 BUFx3_ASAP7_75t_R place2835 (.A(_06376_),
    .Y(net2835));
 BUFx3_ASAP7_75t_R place2833 (.A(net5505),
    .Y(net2833));
 BUFx3_ASAP7_75t_R place2832 (.A(_02344_),
    .Y(net2832));
 BUFx3_ASAP7_75t_R place2831 (.A(_02347_),
    .Y(net2831));
 BUFx3_ASAP7_75t_R place2834 (.A(_06406_),
    .Y(net2834));
 BUFx3_ASAP7_75t_R place2829 (.A(_04045_),
    .Y(net2829));
 BUFx6f_ASAP7_75t_R place2828 (.A(_04053_),
    .Y(net2828));
 BUFx3_ASAP7_75t_R place2827 (.A(net5685),
    .Y(net2827));
 BUFx6f_ASAP7_75t_R place2825 (.A(_06352_),
    .Y(net2825));
 BUFx3_ASAP7_75t_R place2824 (.A(_06374_),
    .Y(net2824));
 BUFx3_ASAP7_75t_R place2822 (.A(_06409_),
    .Y(net2822));
 BUFx3_ASAP7_75t_R place2823 (.A(_06387_),
    .Y(net2823));
 BUFx3_ASAP7_75t_R place2821 (.A(net5431),
    .Y(net2821));
 BUFx3_ASAP7_75t_R place2820 (.A(_02360_),
    .Y(net2820));
 BUFx3_ASAP7_75t_R place2819 (.A(_02361_),
    .Y(net2819));
 BUFx3_ASAP7_75t_R place2817 (.A(_04057_),
    .Y(net2817));
 BUFx3_ASAP7_75t_R place2816 (.A(_04067_),
    .Y(net2816));
 BUFx3_ASAP7_75t_R place2815 (.A(_04081_),
    .Y(net2815));
 BUFx3_ASAP7_75t_R place2814 (.A(_05257_),
    .Y(net2814));
 BUFx3_ASAP7_75t_R place2813 (.A(_05272_),
    .Y(net2813));
 BUFx3_ASAP7_75t_R place2811 (.A(_05297_),
    .Y(net2811));
 BUFx3_ASAP7_75t_R place2810 (.A(net5876),
    .Y(net2810));
 BUFx3_ASAP7_75t_R place2809 (.A(_02369_),
    .Y(net2809));
 BUFx3_ASAP7_75t_R place2808 (.A(_02382_),
    .Y(net2808));
 BUFx3_ASAP7_75t_R place2807 (.A(net5420),
    .Y(net2807));
 BUFx3_ASAP7_75t_R place2806 (.A(_02396_),
    .Y(net2806));
 BUFx3_ASAP7_75t_R place2805 (.A(_04040_),
    .Y(net2805));
 BUFx3_ASAP7_75t_R place2804 (.A(_04062_),
    .Y(net2804));
 BUFx3_ASAP7_75t_R place2803 (.A(_04068_),
    .Y(net2803));
 BUFx3_ASAP7_75t_R place2802 (.A(net5718),
    .Y(net2802));
 BUFx3_ASAP7_75t_R place2800 (.A(_04116_),
    .Y(net2800));
 BUFx3_ASAP7_75t_R place2799 (.A(_05292_),
    .Y(net2799));
 BUFx3_ASAP7_75t_R place2798 (.A(_06404_),
    .Y(net2798));
 BUFx3_ASAP7_75t_R place2797 (.A(_06408_),
    .Y(net2797));
 BUFx3_ASAP7_75t_R place2796 (.A(_02346_),
    .Y(net2796));
 BUFx3_ASAP7_75t_R place2795 (.A(_02358_),
    .Y(net2795));
 BUFx3_ASAP7_75t_R place2794 (.A(_02374_),
    .Y(net2794));
 BUFx3_ASAP7_75t_R place2793 (.A(_02381_),
    .Y(net2793));
 BUFx3_ASAP7_75t_R place2790 (.A(_04071_),
    .Y(net2790));
 BUFx3_ASAP7_75t_R place2789 (.A(_04079_),
    .Y(net2789));
 BUFx3_ASAP7_75t_R place2788 (.A(net5720),
    .Y(net2788));
 BUFx3_ASAP7_75t_R place2786 (.A(_04117_),
    .Y(net2786));
 BUFx3_ASAP7_75t_R place2785 (.A(_05296_),
    .Y(net2785));
 BUFx3_ASAP7_75t_R place2784 (.A(net5964),
    .Y(net2784));
 BUFx3_ASAP7_75t_R place2783 (.A(net5622),
    .Y(net2783));
 BUFx3_ASAP7_75t_R place2782 (.A(_06422_),
    .Y(net2782));
 BUFx3_ASAP7_75t_R place2779 (.A(_04094_),
    .Y(net2779));
 BUFx3_ASAP7_75t_R place2778 (.A(_04118_),
    .Y(net2778));
 BUFx3_ASAP7_75t_R place2777 (.A(_05295_),
    .Y(net2777));
 BUFx3_ASAP7_75t_R place2776 (.A(_05313_),
    .Y(net2776));
 BUFx3_ASAP7_75t_R place2774 (.A(_05318_),
    .Y(net2774));
 BUFx3_ASAP7_75t_R place2773 (.A(_05330_),
    .Y(net2773));
 BUFx3_ASAP7_75t_R place2772 (.A(_05336_),
    .Y(net2772));
 BUFx3_ASAP7_75t_R place2771 (.A(net5598),
    .Y(net2771));
 BUFx3_ASAP7_75t_R place2769 (.A(_06421_),
    .Y(net2769));
 BUFx3_ASAP7_75t_R place2768 (.A(_06434_),
    .Y(net2768));
 BUFx3_ASAP7_75t_R place2770 (.A(_06412_),
    .Y(net2770));
 BUFx6f_ASAP7_75t_R place2767 (.A(_02371_),
    .Y(net2767));
 BUFx6f_ASAP7_75t_R place2765 (.A(_02387_),
    .Y(net2765));
 BUFx3_ASAP7_75t_R place2762 (.A(_04087_),
    .Y(net2762));
 BUFx3_ASAP7_75t_R place2760 (.A(_05314_),
    .Y(net2760));
 BUFx6f_ASAP7_75t_R place2758 (.A(_06423_),
    .Y(net2758));
 BUFx3_ASAP7_75t_R place2756 (.A(net5702),
    .Y(net2756));
 BUFx3_ASAP7_75t_R place2755 (.A(_04106_),
    .Y(net2755));
 BUFx3_ASAP7_75t_R place2754 (.A(_04130_),
    .Y(net2754));
 BUFx3_ASAP7_75t_R place2752 (.A(_04136_),
    .Y(net2752));
 BUFx3_ASAP7_75t_R place2751 (.A(_04192_),
    .Y(net2751));
 BUFx3_ASAP7_75t_R place2750 (.A(_06439_),
    .Y(net2750));
 BUFx3_ASAP7_75t_R place2747 (.A(_04107_),
    .Y(net2747));
 BUFx6f_ASAP7_75t_R rebuffer6028 (.A(net4016),
    .Y(net6028));
 BUFx3_ASAP7_75t_R place2745 (.A(_04131_),
    .Y(net2745));
 BUFx6f_ASAP7_75t_R place2743 (.A(_05319_),
    .Y(net2743));
 BUFx3_ASAP7_75t_R place2742 (.A(_05327_),
    .Y(net2742));
 BUFx3_ASAP7_75t_R place2741 (.A(_06442_),
    .Y(net2741));
 BUFx3_ASAP7_75t_R rebuffer5731 (.A(_02506_),
    .Y(net5731));
 BUFx3_ASAP7_75t_R place2740 (.A(_06451_),
    .Y(net2740));
 BUFx3_ASAP7_75t_R place2739 (.A(_06456_),
    .Y(net2739));
 BUFx3_ASAP7_75t_R place2748 (.A(_06448_),
    .Y(net2748));
 BUFx3_ASAP7_75t_R place2738 (.A(net5693),
    .Y(net2738));
 BUFx3_ASAP7_75t_R place2736 (.A(_05340_),
    .Y(net2736));
 BUFx3_ASAP7_75t_R place2737 (.A(_05329_),
    .Y(net2737));
 BUFx3_ASAP7_75t_R place2733 (.A(_06453_),
    .Y(net2733));
 BUFx3_ASAP7_75t_R place2732 (.A(_04142_),
    .Y(net2732));
 BUFx3_ASAP7_75t_R place2731 (.A(_05325_),
    .Y(net2731));
 BUFx3_ASAP7_75t_R place2730 (.A(_05342_),
    .Y(net2730));
 BUFx3_ASAP7_75t_R place2729 (.A(_05361_),
    .Y(net2729));
 BUFx3_ASAP7_75t_R rebuffer5725 (.A(net2764),
    .Y(net5725));
 BUFx3_ASAP7_75t_R place2727 (.A(_06461_),
    .Y(net2727));
 BUFx3_ASAP7_75t_R rebuffer5730 (.A(_00529_),
    .Y(net5730));
 BUFx3_ASAP7_75t_R place2735 (.A(net2734),
    .Y(net2735));
 BUFx3_ASAP7_75t_R place2734 (.A(_05346_),
    .Y(net2734));
 BUFx3_ASAP7_75t_R place2725 (.A(_02492_),
    .Y(net2725));
 BUFx6f_ASAP7_75t_R place2723 (.A(_04143_),
    .Y(net2723));
 BUFx3_ASAP7_75t_R place2722 (.A(_05343_),
    .Y(net2722));
 BUFx3_ASAP7_75t_R place2720 (.A(_05360_),
    .Y(net2720));
 BUFx3_ASAP7_75t_R place2719 (.A(_05365_),
    .Y(net2719));
 BUFx3_ASAP7_75t_R place2718 (.A(_02522_),
    .Y(net2718));
 BUFx6f_ASAP7_75t_R place2724 (.A(_04143_),
    .Y(net2724));
 BUFx3_ASAP7_75t_R place2721 (.A(_05348_),
    .Y(net2721));
 BUFx6f_ASAP7_75t_R place2715 (.A(_06470_),
    .Y(net2715));
 BUFx6f_ASAP7_75t_R place2714 (.A(_06470_),
    .Y(net2714));
 BUFx3_ASAP7_75t_R rebuffer6027 (.A(_02895_),
    .Y(net6027));
 BUFx12f_ASAP7_75t_R place2711 (.A(net5419),
    .Y(net2711));
 BUFx3_ASAP7_75t_R place2712 (.A(net5419),
    .Y(net2712));
 BUFx6f_ASAP7_75t_R place2709 (.A(_04329_),
    .Y(net2709));
 BUFx6f_ASAP7_75t_R place2708 (.A(_04125_),
    .Y(net2708));
 BUFx6f_ASAP7_75t_R place2707 (.A(_04125_),
    .Y(net2707));
 BUFx3_ASAP7_75t_R place2706 (.A(_05370_),
    .Y(net2706));
 BUFx6f_ASAP7_75t_R place2704 (.A(_02524_),
    .Y(net2704));
 BUFx12f_ASAP7_75t_R place2713 (.A(net5372),
    .Y(net2713));
 BUFx12f_ASAP7_75t_R place2710 (.A(net5592),
    .Y(net2710));
 BUFx6f_ASAP7_75t_R place2703 (.A(_03065_),
    .Y(net2703));
 BUFx12f_ASAP7_75t_R place2705 (.A(_02524_),
    .Y(net2705));
 BUFx12f_ASAP7_75t_R place2699 (.A(_04330_),
    .Y(net2699));
 BUFx6f_ASAP7_75t_R place2697 (.A(_05374_),
    .Y(net2697));
 BUFx12f_ASAP7_75t_R place2700 (.A(_04330_),
    .Y(net2700));
 BUFx6f_ASAP7_75t_R place2698 (.A(_05374_),
    .Y(net2698));
 BUFx6f_ASAP7_75t_R place2696 (.A(_05355_),
    .Y(net2696));
 BUFx12f_ASAP7_75t_R place2702 (.A(_04330_),
    .Y(net2702));
 BUFx24_ASAP7_75t_R clkbuf_leaf_1_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_1_clk));
 BUFx3_ASAP7_75t_R place2701 (.A(net5910),
    .Y(net2701));
 BUFx24_ASAP7_75t_R clkbuf_leaf_0_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_0_clk));
 BUFx6f_ASAP7_75t_R place2717 (.A(_06457_),
    .Y(net2717));
 BUFx6f_ASAP7_75t_R place2716 (.A(_06457_),
    .Y(net2716));
 BUFx2_ASAP7_75t_R output213 (.A(net213),
    .Y(mfcc_done_o));
 BUFx2_ASAP7_75t_R input212 (.A(start_i),
    .Y(net212));
 BUFx2_ASAP7_75t_R input211 (.A(rst_n),
    .Y(net211));
 BUFx2_ASAP7_75t_R input210 (.A(pcm_ready_i),
    .Y(net210));
 BUFx2_ASAP7_75t_R input209 (.A(auto_restart_i),
    .Y(net209));
 DFFHQNx1_ASAP7_75t_R \hamming_finished$_SDFFE_PP0P_  (.CLK(clknet_leaf_20_clk),
    .D(_00557_),
    .QN(_00317_));
 DFFHQNx1_ASAP7_75t_R \start_move$_DFFE_PN_  (.CLK(clknet_leaf_20_clk),
    .D(_00558_),
    .QN(_00316_));
 DFFHQNx1_ASAP7_75t_R \start_move_auto$_SDFF_PN0_  (.CLK(clknet_leaf_18_clk),
    .D(_00559_),
    .QN(_00315_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.read_ptr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00560_),
    .QN(_00543_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.read_ptr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_00561_),
    .QN(_00544_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.read_ptr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00562_),
    .QN(_00314_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.read_ptr[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00563_),
    .QN(_00313_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.read_ptr[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00564_),
    .QN(_00312_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.read_ptr[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00565_),
    .QN(_00311_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.read_ptr[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00566_),
    .QN(_00310_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.read_ptr[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_00567_),
    .QN(_00309_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.write_ptr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00568_),
    .QN(_00069_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.write_ptr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_00569_),
    .QN(_00308_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.write_ptr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00570_),
    .QN(_00307_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.write_ptr[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00571_),
    .QN(_00306_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.write_ptr[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00572_),
    .QN(_00305_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.write_ptr[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_00573_),
    .QN(_00304_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.write_ptr[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_00574_),
    .QN(_00303_));
 DFFHQNx1_ASAP7_75t_R \tx_fifo.write_ptr[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_00575_),
    .QN(_00302_));
 DFFHQNx1_ASAP7_75t_R \u_dct.dct_done_o$_SDFF_PN0_  (.CLK(clknet_leaf_6_clk),
    .D(_00576_),
    .QN(_00318_));
 DFFHQNx1_ASAP7_75t_R \u_dct.dct_state[0]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00006_),
    .QN(_00319_));
 DFFHQNx1_ASAP7_75t_R \u_dct.dct_state[1]$_DFF_P_  (.CLK(clknet_leaf_9_clk),
    .D(_00000_),
    .QN(_00320_));
 DFFHQNx1_ASAP7_75t_R \u_dct.dct_state[2]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00007_),
    .QN(_00321_));
 DFFHQNx1_ASAP7_75t_R \u_dct.dct_state[3]$_DFF_P_  (.CLK(clknet_leaf_7_clk),
    .D(_00001_),
    .QN(_00301_));
 DFFHQNx1_ASAP7_75t_R \u_dct.k_ptr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_00577_),
    .QN(_00470_));
 DFFHQNx1_ASAP7_75t_R \u_dct.k_ptr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_00578_),
    .QN(_00471_));
 DFFHQNx1_ASAP7_75t_R \u_dct.k_ptr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_00579_),
    .QN(_00300_));
 DFFHQNx1_ASAP7_75t_R \u_dct.k_ptr[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_00580_),
    .QN(_00299_));
 DFFHQNx1_ASAP7_75t_R \u_dct.n_ptr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_00581_),
    .QN(_00475_));
 DFFHQNx1_ASAP7_75t_R \u_dct.n_ptr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_00582_),
    .QN(_00476_));
 DFFHQNx1_ASAP7_75t_R \u_dct.n_ptr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_00583_),
    .QN(_00298_));
 DFFHQNx1_ASAP7_75t_R \u_dct.n_ptr[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_00584_),
    .QN(_00297_));
 DFFHQNx1_ASAP7_75t_R \u_dct.n_ptr[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_00585_),
    .QN(_00296_));
 DFFHQNx1_ASAP7_75t_R \u_dct.n_ptr[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_00586_),
    .QN(_00295_));
 DFFHQNx1_ASAP7_75t_R \u_fft.fft_done_o$_SDFF_PN0_  (.CLK(clknet_leaf_5_clk),
    .D(_00587_),
    .QN(_00322_));
 DFFHQNx1_ASAP7_75t_R \u_fft.fft_state[0]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00008_),
    .QN(_00323_));
 DFFHQNx1_ASAP7_75t_R \u_fft.fft_state[1]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00009_),
    .QN(_00324_));
 DFFHQNx1_ASAP7_75t_R \u_fft.fft_state[2]$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(_00010_),
    .QN(_00068_));
 DFFHQNx1_ASAP7_75t_R \u_fft.fft_state[3]$_DFF_P_  (.CLK(clknet_leaf_1_clk),
    .D(_00002_),
    .QN(_00294_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_00588_),
    .QN(_00293_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00589_),
    .QN(_00292_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00590_),
    .QN(_00291_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_00591_),
    .QN(_00290_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .D(_00592_),
    .QN(_00289_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_00593_),
    .QN(_00288_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_00594_),
    .QN(_00287_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_00595_),
    .QN(_00286_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_00596_),
    .QN(_00285_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_00597_),
    .QN(_00284_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage1[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_00598_),
    .QN(_00283_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage1[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00599_),
    .QN(_00282_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage1[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00600_),
    .QN(_00281_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage1[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_00601_),
    .QN(_00280_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage1[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00602_),
    .QN(_00279_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage1[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_00603_),
    .QN(_00278_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage1[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_00604_),
    .QN(_00277_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage1[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_00605_),
    .QN(_00276_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage1[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_00606_),
    .QN(_00275_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage1[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_5_clk),
    .D(_00607_),
    .QN(_00274_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage2[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00608_),
    .QN(_00273_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage2[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00609_),
    .QN(_00272_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage2[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00610_),
    .QN(_00271_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage2[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_00611_),
    .QN(_00270_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage2[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00612_),
    .QN(_00269_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage2[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00613_),
    .QN(_00268_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage2[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00614_),
    .QN(_00267_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage2[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00615_),
    .QN(_00266_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage2[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00616_),
    .QN(_00265_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage2[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00617_),
    .QN(_00264_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage3[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00618_),
    .QN(_00263_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage3[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00619_),
    .QN(_00262_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage3[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00620_),
    .QN(_00261_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage3[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_00621_),
    .QN(_00260_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage3[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00622_),
    .QN(_00259_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage3[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00623_),
    .QN(_00258_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage3[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00624_),
    .QN(_00257_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage3[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00625_),
    .QN(_00256_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage3[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00626_),
    .QN(_00255_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage3[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00627_),
    .QN(_00254_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage4[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00628_),
    .QN(_00253_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage4[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00629_),
    .QN(_00252_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage4[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00630_),
    .QN(_00251_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage4[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00631_),
    .QN(_00250_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage4[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00632_),
    .QN(_00249_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage4[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00633_),
    .QN(_00248_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage4[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_00634_),
    .QN(_00247_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage4[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00635_),
    .QN(_00246_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage4[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00636_),
    .QN(_00245_));
 DFFHQNx1_ASAP7_75t_R \u_fft.power_ptr_stage4[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .D(_00637_),
    .QN(_00244_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[20]$_SDFFE_PN1P_  (.CLK(clknet_leaf_26_clk),
    .D(_00638_),
    .QN(_00365_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_00639_),
    .QN(_00366_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_00640_),
    .QN(_00243_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_00641_),
    .QN(_00242_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_00642_),
    .QN(_00241_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_00643_),
    .QN(_00240_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_00644_),
    .QN(_00239_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_00645_),
    .QN(_00238_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_00646_),
    .QN(_00237_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_00647_),
    .QN(_00236_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_00648_),
    .QN(_00396_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[31]$_SDFFE_PN1P_  (.CLK(clknet_leaf_0_clk),
    .D(_00649_),
    .QN(_00397_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[32]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_00650_),
    .QN(_00235_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[33]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_00651_),
    .QN(_00234_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[34]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_00652_),
    .QN(_00233_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[35]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_00653_),
    .QN(_00232_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[36]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_00654_),
    .QN(_00231_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[37]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_00655_),
    .QN(_00230_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[38]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_00656_),
    .QN(_00229_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[39]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_00657_),
    .QN(_00228_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[40]$_SDFFE_PN1P_  (.CLK(clknet_leaf_27_clk),
    .D(_00658_),
    .QN(_00480_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[41]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_00659_),
    .QN(_00481_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[42]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_00660_),
    .QN(_00488_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[43]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_00661_),
    .QN(_00057_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[44]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_00662_),
    .QN(_00067_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[45]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_00663_),
    .QN(_00227_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[46]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_00664_),
    .QN(_00226_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[47]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_00665_),
    .QN(_00066_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[48]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_00666_),
    .QN(_00225_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[49]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_00667_),
    .QN(_00065_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[50]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_00668_),
    .QN(_00064_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[51]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_00669_),
    .QN(_00063_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[52]$_SDFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_00670_),
    .QN(_00224_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[53]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_00671_),
    .QN(_00062_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[54]$_SDFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .D(_00672_),
    .QN(_00061_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[55]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_00673_),
    .QN(_00494_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[56]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_00674_),
    .QN(_00223_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[57]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_00675_),
    .QN(_00222_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[58]$_SDFFE_PN0P_  (.CLK(clknet_leaf_0_clk),
    .D(_00676_),
    .QN(_00221_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[59]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_00677_),
    .QN(_00220_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[60]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_00678_),
    .QN(_00219_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[61]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_00679_),
    .QN(_00218_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[62]$_SDFFE_PN0P_  (.CLK(clknet_leaf_1_clk),
    .D(_00680_),
    .QN(_00217_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[63]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_00681_),
    .QN(_00216_));
 DFFHQNx1_ASAP7_75t_R \u_fft.sched[64]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_00682_),
    .QN(_00215_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00683_),
    .QN(_00548_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[10]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00684_),
    .QN(_00214_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[11]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00685_),
    .QN(_00213_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[12]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_00686_),
    .QN(_00212_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[13]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00687_),
    .QN(_00211_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[14]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00688_),
    .QN(_00210_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[15]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_00689_),
    .QN(_00209_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[16]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00690_),
    .QN(_00208_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[17]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_00691_),
    .QN(_00207_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[18]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .D(_00692_),
    .QN(_00206_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[19]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00693_),
    .QN(_00205_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00694_),
    .QN(_00549_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[20]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00695_),
    .QN(_00204_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[21]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00696_),
    .QN(_00203_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[22]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00697_),
    .QN(_00202_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[23]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00698_),
    .QN(_00201_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[24]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00699_),
    .QN(_00200_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[25]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00700_),
    .QN(_00199_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[26]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00701_),
    .QN(_00198_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[27]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00702_),
    .QN(_00197_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[28]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00703_),
    .QN(_00196_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[29]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00704_),
    .QN(_00195_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_00705_),
    .QN(_00194_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[30]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .D(_00706_),
    .QN(_00193_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[31]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00707_),
    .QN(_00192_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00708_),
    .QN(_00191_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00709_),
    .QN(_00190_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00710_),
    .QN(_00189_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00711_),
    .QN(_00188_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00712_),
    .QN(_00187_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[8]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00713_),
    .QN(_00186_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.calc_pointer[9]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00714_),
    .QN(_00185_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.done$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .D(_00715_),
    .QN(_00325_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.done_o$_DFF_P_  (.CLK(clknet_leaf_2_clk),
    .D(\u_hamming_window.done ),
    .QN(_00184_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.frame_ptr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_00716_),
    .QN(_00024_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.frame_ptr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_00717_),
    .QN(_00183_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.frame_ptr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00718_),
    .QN(_00182_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.frame_ptr[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .D(_00719_),
    .QN(_00181_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.frame_ptr[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .D(_00720_),
    .QN(_00180_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.frame_ptr[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_00721_),
    .QN(_00179_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.frame_ptr[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .D(_00722_),
    .QN(_00178_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.frame_ptr[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_00723_),
    .QN(_00177_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.frame_ptr[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_00724_),
    .QN(_00326_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.hamming_state[0]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00011_),
    .QN(_00327_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.hamming_state[1]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00012_),
    .QN(_00328_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.hamming_state[2]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00013_),
    .QN(_00046_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.hamming_state[3]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .D(_00003_),
    .QN(_00176_));
 DFFHQNx1_ASAP7_75t_R \u_hamming_window.rd_en_o$_SDFF_PN0_  (.CLK(clknet_leaf_20_clk),
    .D(_00725_),
    .QN(_00175_));
 DFFHQNx1_ASAP7_75t_R \u_mel.k[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_00726_),
    .QN(\u_mel.k_next[0] ));
 DFFHQNx1_ASAP7_75t_R \u_mel.k[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .D(_00727_),
    .QN(_00553_));
 DFFHQNx1_ASAP7_75t_R \u_mel.k[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_00728_),
    .QN(_00174_));
 DFFHQNx1_ASAP7_75t_R \u_mel.k[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_00729_),
    .QN(_00173_));
 DFFHQNx1_ASAP7_75t_R \u_mel.k[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_00730_),
    .QN(_00172_));
 DFFHQNx1_ASAP7_75t_R \u_mel.k[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_00731_),
    .QN(_00171_));
 DFFHQNx1_ASAP7_75t_R \u_mel.k[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_00732_),
    .QN(_00170_));
 DFFHQNx1_ASAP7_75t_R \u_mel.k[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .D(_00733_),
    .QN(_00169_));
 DFFHQNx1_ASAP7_75t_R \u_mel.k[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_00734_),
    .QN(_00168_));
 DFFHQNx1_ASAP7_75t_R \u_mel.mel_done_o$_SDFF_PN0_  (.CLK(clknet_leaf_7_clk),
    .D(_00735_),
    .QN(_00167_));
 DFFHQNx1_ASAP7_75t_R \u_mel.mel_prt_energies[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_00736_),
    .QN(_00518_));
 DFFHQNx1_ASAP7_75t_R \u_mel.mel_prt_energies[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_00737_),
    .QN(_00519_));
 DFFHQNx1_ASAP7_75t_R \u_mel.mel_prt_energies[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_00738_),
    .QN(_00166_));
 DFFHQNx1_ASAP7_75t_R \u_mel.mel_prt_energies[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_00739_),
    .QN(_00165_));
 DFFHQNx1_ASAP7_75t_R \u_mel.mel_prt_energies[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .D(_00740_),
    .QN(_00164_));
 DFFHQNx1_ASAP7_75t_R \u_mel.mel_prt_energies[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .D(_00741_),
    .QN(_00329_));
 DFFHQNx1_ASAP7_75t_R \u_mel.state[0]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00014_),
    .QN(_00330_));
 DFFHQNx1_ASAP7_75t_R \u_mel.state[1]$_DFF_P_  (.CLK(clknet_leaf_8_clk),
    .D(_00015_),
    .QN(_00331_));
 DFFHQNx1_ASAP7_75t_R \u_mel.state[2]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00016_),
    .QN(_00332_));
 DFFHQNx1_ASAP7_75t_R \u_mel.state[3]$_DFF_P_  (.CLK(clknet_leaf_5_clk),
    .D(_00004_),
    .QN(_00163_));
 DFFHQNx1_ASAP7_75t_R \u_pre_emphasis.out_valid$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .D(_00742_),
    .QN(_00333_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.current_state[0]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(net5360),
    .QN(_00334_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.current_state[1]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00018_),
    .QN(_00335_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.current_state[2]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00019_),
    .QN(_00055_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.current_state[3]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(_00005_),
    .QN(_00336_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.current_state[4]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .D(net4374),
    .QN(_00162_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.fifo_rd_en_o$_SDFF_PN0_  (.CLK(clknet_leaf_2_clk),
    .D(_00743_),
    .QN(_00161_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[10]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00744_),
    .QN(_00160_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[11]$_SDFFE_PN0N_  (.CLK(clknet_leaf_15_clk),
    .D(_00745_),
    .QN(_00159_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[12]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00746_),
    .QN(_00158_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[13]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00747_),
    .QN(_00157_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[14]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00748_),
    .QN(_00156_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[15]$_SDFFE_PN0N_  (.CLK(clknet_leaf_15_clk),
    .D(_00749_),
    .QN(_00155_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[16]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00750_),
    .QN(_00154_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[17]$_SDFFE_PN0N_  (.CLK(clknet_leaf_15_clk),
    .D(_00751_),
    .QN(_00153_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[18]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00752_),
    .QN(_00152_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[19]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00753_),
    .QN(_00151_));
 DFFHQNx2_ASAP7_75t_R \u_window_buffer.internal_read_ptr[1]$_SDFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .D(_00754_),
    .QN(_00523_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[20]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00755_),
    .QN(_00150_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[21]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00756_),
    .QN(_00149_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[22]$_SDFFE_PN0N_  (.CLK(clknet_leaf_12_clk),
    .D(_00757_),
    .QN(_00148_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[23]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00758_),
    .QN(_00147_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[24]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00759_),
    .QN(_00146_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[25]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00760_),
    .QN(_00145_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[26]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00761_),
    .QN(_00144_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[27]$_SDFFE_PN0N_  (.CLK(clknet_leaf_13_clk),
    .D(_00762_),
    .QN(_00143_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[28]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00763_),
    .QN(_00142_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[29]$_SDFFE_PN0N_  (.CLK(clknet_leaf_13_clk),
    .D(_00764_),
    .QN(_00141_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[2]$_SDFFE_PN0N_  (.CLK(clknet_leaf_15_clk),
    .D(_00765_),
    .QN(_00524_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[30]$_SDFFE_PN0N_  (.CLK(clknet_leaf_13_clk),
    .D(_00766_),
    .QN(_00140_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[31]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00767_),
    .QN(_00139_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[3]$_SDFFE_PN0N_  (.CLK(clknet_leaf_15_clk),
    .D(_00768_),
    .QN(_00058_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[4]$_SDFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .D(_00769_),
    .QN(_00059_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[5]$_SDFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .D(_00770_),
    .QN(_00138_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[6]$_SDFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .D(_00771_),
    .QN(_00137_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[7]$_SDFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .D(_00772_),
    .QN(_00136_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[8]$_SDFFE_PN0N_  (.CLK(clknet_leaf_10_clk),
    .D(_00773_),
    .QN(_00135_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.internal_read_ptr[9]$_SDFFE_PN0N_  (.CLK(clknet_leaf_14_clk),
    .D(_00774_),
    .QN(_00134_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_00775_),
    .QN(_00534_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_00776_),
    .QN(_00133_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_00777_),
    .QN(_00132_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00778_),
    .QN(_00131_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00779_),
    .QN(_00130_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_00780_),
    .QN(_00129_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00781_),
    .QN(_00128_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00782_),
    .QN(_00127_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00783_),
    .QN(_00126_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00784_),
    .QN(_00125_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00785_),
    .QN(_00124_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_00786_),
    .QN(_00535_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00787_),
    .QN(_00123_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00788_),
    .QN(_00122_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_00789_),
    .QN(_00121_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_00790_),
    .QN(_00120_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00791_),
    .QN(_00119_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_00792_),
    .QN(_00118_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_00793_),
    .QN(_00117_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_00794_),
    .QN(_00116_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .D(_00795_),
    .QN(_00115_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_00796_),
    .QN(_00114_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_00797_),
    .QN(_00113_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_00798_),
    .QN(_00112_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .D(_00799_),
    .QN(_00111_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_00800_),
    .QN(_00110_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_00801_),
    .QN(_00109_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_00802_),
    .QN(_00108_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_00803_),
    .QN(_00107_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_00804_),
    .QN(_00106_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_00805_),
    .QN(_00105_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.move_counter[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .D(_00806_),
    .QN(_00337_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.next_state_is_valid_to_read$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .D(_00023_),
    .QN(_00104_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_00807_),
    .QN(_00461_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_00808_),
    .QN(_00103_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_00809_),
    .QN(_00102_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_00810_),
    .QN(_00101_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_00811_),
    .QN(_00100_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_00812_),
    .QN(_00099_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_00813_),
    .QN(_00098_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_00814_),
    .QN(_00097_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_00815_),
    .QN(_00096_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_00816_),
    .QN(_00095_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_00817_),
    .QN(_00094_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_00818_),
    .QN(_00093_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_00819_),
    .QN(_00092_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_00820_),
    .QN(_00091_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_00821_),
    .QN(_00090_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_00822_),
    .QN(_00089_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_00823_),
    .QN(_00088_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_00824_),
    .QN(_00087_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_00825_),
    .QN(_00086_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .D(_00826_),
    .QN(_00085_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .D(_00827_),
    .QN(_00084_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .D(_00828_),
    .QN(_00083_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_00829_),
    .QN(_00082_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .D(_00830_),
    .QN(_00081_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .D(_00831_),
    .QN(_00080_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .D(_00832_),
    .QN(_00079_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_00833_),
    .QN(_00078_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_00834_),
    .QN(_00077_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_00835_),
    .QN(_00076_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_00836_),
    .QN(_00075_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_00837_),
    .QN(_00074_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.read_ptr[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .D(_00838_),
    .QN(_00073_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.start_next_state_o$_SDFF_PN0_  (.CLK(clknet_leaf_21_clk),
    .D(_00839_),
    .QN(_00072_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_00840_),
    .QN(_00872_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_00841_),
    .QN(_00031_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_00842_),
    .QN(_00032_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_00843_),
    .QN(_00033_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_00844_),
    .QN(_00034_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_00845_),
    .QN(_00035_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_00846_),
    .QN(_00036_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_00847_),
    .QN(_00037_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_00848_),
    .QN(_00038_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_00849_),
    .QN(_00039_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_00850_),
    .QN(_00040_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_00851_),
    .QN(_00071_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_00852_),
    .QN(_00041_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_00853_),
    .QN(_00042_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_00854_),
    .QN(_00043_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_00855_),
    .QN(_00044_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_00856_),
    .QN(_00045_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_00857_),
    .QN(_00047_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_00858_),
    .QN(_00048_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_00859_),
    .QN(_00049_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .D(_00860_),
    .QN(_00050_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_00861_),
    .QN(_00051_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_00862_),
    .QN(_00060_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .D(_00863_),
    .QN(_00052_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_00864_),
    .QN(_00053_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_00865_),
    .QN(_00070_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_00866_),
    .QN(_00025_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_00867_),
    .QN(_00026_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_00868_),
    .QN(_00027_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_16_clk),
    .D(_00869_),
    .QN(_00028_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_00870_),
    .QN(_00029_));
 DFFHQNx1_ASAP7_75t_R \u_window_buffer.write_ptr[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_17_clk),
    .D(_00871_),
    .QN(_00030_));
 TIELOx1_ASAP7_75t_R _12776__1 (.L(mfcc_data_o[0]));
 TIELOx1_ASAP7_75t_R _12777__2 (.L(mfcc_data_o[1]));
 TIELOx1_ASAP7_75t_R _12778__3 (.L(mfcc_data_o[2]));
 TIELOx1_ASAP7_75t_R _12779__4 (.L(mfcc_data_o[3]));
 TIELOx1_ASAP7_75t_R _12780__5 (.L(mfcc_data_o[4]));
 TIELOx1_ASAP7_75t_R _12781__6 (.L(mfcc_data_o[5]));
 TIELOx1_ASAP7_75t_R _12782__7 (.L(mfcc_data_o[6]));
 TIELOx1_ASAP7_75t_R _12783__8 (.L(mfcc_data_o[7]));
 TIELOx1_ASAP7_75t_R _12784__9 (.L(mfcc_data_o[8]));
 TIELOx1_ASAP7_75t_R _12785__10 (.L(mfcc_data_o[9]));
 TIELOx1_ASAP7_75t_R _12786__11 (.L(mfcc_data_o[10]));
 TIELOx1_ASAP7_75t_R _12787__12 (.L(mfcc_data_o[11]));
 TIELOx1_ASAP7_75t_R _12788__13 (.L(mfcc_data_o[12]));
 TIELOx1_ASAP7_75t_R _12789__14 (.L(mfcc_data_o[13]));
 TIELOx1_ASAP7_75t_R _12790__15 (.L(mfcc_data_o[14]));
 TIELOx1_ASAP7_75t_R _12791__16 (.L(mfcc_data_o[15]));
 TIELOx1_ASAP7_75t_R _12792__17 (.L(mfcc_data_o[16]));
 TIELOx1_ASAP7_75t_R _12793__18 (.L(mfcc_data_o[17]));
 TIELOx1_ASAP7_75t_R _12794__19 (.L(mfcc_data_o[18]));
 TIELOx1_ASAP7_75t_R _12795__20 (.L(mfcc_data_o[19]));
 TIELOx1_ASAP7_75t_R _12796__21 (.L(mfcc_data_o[20]));
 TIELOx1_ASAP7_75t_R _12797__22 (.L(mfcc_data_o[21]));
 TIELOx1_ASAP7_75t_R _12798__23 (.L(mfcc_data_o[22]));
 TIELOx1_ASAP7_75t_R _12799__24 (.L(mfcc_data_o[23]));
 TIELOx1_ASAP7_75t_R _12800__25 (.L(mfcc_data_o[24]));
 TIELOx1_ASAP7_75t_R _12801__26 (.L(mfcc_data_o[25]));
 TIELOx1_ASAP7_75t_R _12802__27 (.L(mfcc_data_o[26]));
 TIELOx1_ASAP7_75t_R _12803__28 (.L(mfcc_data_o[27]));
 TIELOx1_ASAP7_75t_R _12804__29 (.L(mfcc_data_o[28]));
 TIELOx1_ASAP7_75t_R _12805__30 (.L(mfcc_data_o[29]));
 TIELOx1_ASAP7_75t_R _12806__31 (.L(mfcc_data_o[30]));
 TIELOx1_ASAP7_75t_R _12807__32 (.L(mfcc_data_o[31]));
 TIELOx1_ASAP7_75t_R _12808__33 (.L(mfcc_data_o[32]));
 TIELOx1_ASAP7_75t_R _12809__34 (.L(mfcc_data_o[33]));
 TIELOx1_ASAP7_75t_R _12810__35 (.L(mfcc_data_o[34]));
 TIELOx1_ASAP7_75t_R _12811__36 (.L(mfcc_data_o[35]));
 TIELOx1_ASAP7_75t_R _12812__37 (.L(mfcc_data_o[36]));
 TIELOx1_ASAP7_75t_R _12813__38 (.L(mfcc_data_o[37]));
 TIELOx1_ASAP7_75t_R _12814__39 (.L(mfcc_data_o[38]));
 TIELOx1_ASAP7_75t_R _12815__40 (.L(mfcc_data_o[39]));
 TIELOx1_ASAP7_75t_R _12816__41 (.L(mfcc_data_o[40]));
 TIELOx1_ASAP7_75t_R _12817__42 (.L(mfcc_data_o[41]));
 TIELOx1_ASAP7_75t_R _12818__43 (.L(mfcc_data_o[42]));
 TIELOx1_ASAP7_75t_R _12819__44 (.L(mfcc_data_o[43]));
 TIELOx1_ASAP7_75t_R _12820__45 (.L(mfcc_data_o[44]));
 TIELOx1_ASAP7_75t_R _12821__46 (.L(mfcc_data_o[45]));
 TIELOx1_ASAP7_75t_R _12822__47 (.L(mfcc_data_o[46]));
 TIELOx1_ASAP7_75t_R _12823__48 (.L(mfcc_data_o[47]));
 TIELOx1_ASAP7_75t_R _12824__49 (.L(mfcc_data_o[48]));
 TIELOx1_ASAP7_75t_R _12825__50 (.L(mfcc_data_o[49]));
 TIELOx1_ASAP7_75t_R _12826__51 (.L(mfcc_data_o[50]));
 TIELOx1_ASAP7_75t_R _12827__52 (.L(mfcc_data_o[51]));
 TIELOx1_ASAP7_75t_R _12828__53 (.L(mfcc_data_o[52]));
 TIELOx1_ASAP7_75t_R _12829__54 (.L(mfcc_data_o[53]));
 TIELOx1_ASAP7_75t_R _12830__55 (.L(mfcc_data_o[54]));
 TIELOx1_ASAP7_75t_R _12831__56 (.L(mfcc_data_o[55]));
 TIELOx1_ASAP7_75t_R _12832__57 (.L(mfcc_data_o[56]));
 TIELOx1_ASAP7_75t_R _12833__58 (.L(mfcc_data_o[57]));
 TIELOx1_ASAP7_75t_R _12834__59 (.L(mfcc_data_o[58]));
 TIELOx1_ASAP7_75t_R _12835__60 (.L(mfcc_data_o[59]));
 TIELOx1_ASAP7_75t_R _12836__61 (.L(mfcc_data_o[60]));
 TIELOx1_ASAP7_75t_R _12837__62 (.L(mfcc_data_o[61]));
 TIELOx1_ASAP7_75t_R _12838__63 (.L(mfcc_data_o[62]));
 TIELOx1_ASAP7_75t_R _12839__64 (.L(mfcc_data_o[63]));
 TIELOx1_ASAP7_75t_R _12840__65 (.L(mfcc_data_o[64]));
 TIELOx1_ASAP7_75t_R _12841__66 (.L(mfcc_data_o[65]));
 TIELOx1_ASAP7_75t_R _12842__67 (.L(mfcc_data_o[66]));
 TIELOx1_ASAP7_75t_R _12843__68 (.L(mfcc_data_o[67]));
 TIELOx1_ASAP7_75t_R _12844__69 (.L(mfcc_data_o[68]));
 TIELOx1_ASAP7_75t_R _12845__70 (.L(mfcc_data_o[69]));
 TIELOx1_ASAP7_75t_R _12846__71 (.L(mfcc_data_o[70]));
 TIELOx1_ASAP7_75t_R _12847__72 (.L(mfcc_data_o[71]));
 TIELOx1_ASAP7_75t_R _12848__73 (.L(mfcc_data_o[72]));
 TIELOx1_ASAP7_75t_R _12849__74 (.L(mfcc_data_o[73]));
 TIELOx1_ASAP7_75t_R _12850__75 (.L(mfcc_data_o[74]));
 TIELOx1_ASAP7_75t_R _12851__76 (.L(mfcc_data_o[75]));
 TIELOx1_ASAP7_75t_R _12852__77 (.L(mfcc_data_o[76]));
 TIELOx1_ASAP7_75t_R _12853__78 (.L(mfcc_data_o[77]));
 TIELOx1_ASAP7_75t_R _12854__79 (.L(mfcc_data_o[78]));
 TIELOx1_ASAP7_75t_R _12855__80 (.L(mfcc_data_o[79]));
 TIELOx1_ASAP7_75t_R _12856__81 (.L(mfcc_data_o[80]));
 TIELOx1_ASAP7_75t_R _12857__82 (.L(mfcc_data_o[81]));
 TIELOx1_ASAP7_75t_R _12858__83 (.L(mfcc_data_o[82]));
 TIELOx1_ASAP7_75t_R _12859__84 (.L(mfcc_data_o[83]));
 TIELOx1_ASAP7_75t_R _12860__85 (.L(mfcc_data_o[84]));
 TIELOx1_ASAP7_75t_R _12861__86 (.L(mfcc_data_o[85]));
 TIELOx1_ASAP7_75t_R _12862__87 (.L(mfcc_data_o[86]));
 TIELOx1_ASAP7_75t_R _12863__88 (.L(mfcc_data_o[87]));
 TIELOx1_ASAP7_75t_R _12864__89 (.L(mfcc_data_o[88]));
 TIELOx1_ASAP7_75t_R _12865__90 (.L(mfcc_data_o[89]));
 TIELOx1_ASAP7_75t_R _12866__91 (.L(mfcc_data_o[90]));
 TIELOx1_ASAP7_75t_R _12867__92 (.L(mfcc_data_o[91]));
 TIELOx1_ASAP7_75t_R _12868__93 (.L(mfcc_data_o[92]));
 TIELOx1_ASAP7_75t_R _12869__94 (.L(mfcc_data_o[93]));
 TIELOx1_ASAP7_75t_R _12870__95 (.L(mfcc_data_o[94]));
 TIELOx1_ASAP7_75t_R _12871__96 (.L(mfcc_data_o[95]));
 TIELOx1_ASAP7_75t_R _12872__97 (.L(mfcc_data_o[96]));
 TIELOx1_ASAP7_75t_R _12873__98 (.L(mfcc_data_o[97]));
 TIELOx1_ASAP7_75t_R _12874__99 (.L(mfcc_data_o[98]));
 TIELOx1_ASAP7_75t_R _12875__100 (.L(mfcc_data_o[99]));
 TIELOx1_ASAP7_75t_R _12876__101 (.L(mfcc_data_o[100]));
 TIELOx1_ASAP7_75t_R _12877__102 (.L(mfcc_data_o[101]));
 TIELOx1_ASAP7_75t_R _12878__103 (.L(mfcc_data_o[102]));
 TIELOx1_ASAP7_75t_R _12879__104 (.L(mfcc_data_o[103]));
 TIELOx1_ASAP7_75t_R _12880__105 (.L(mfcc_data_o[104]));
 TIELOx1_ASAP7_75t_R _12881__106 (.L(mfcc_data_o[105]));
 TIELOx1_ASAP7_75t_R _12882__107 (.L(mfcc_data_o[106]));
 TIELOx1_ASAP7_75t_R _12883__108 (.L(mfcc_data_o[107]));
 TIELOx1_ASAP7_75t_R _12884__109 (.L(mfcc_data_o[108]));
 TIELOx1_ASAP7_75t_R _12885__110 (.L(mfcc_data_o[109]));
 TIELOx1_ASAP7_75t_R _12886__111 (.L(mfcc_data_o[110]));
 TIELOx1_ASAP7_75t_R _12887__112 (.L(mfcc_data_o[111]));
 TIELOx1_ASAP7_75t_R _12888__113 (.L(mfcc_data_o[112]));
 TIELOx1_ASAP7_75t_R _12889__114 (.L(mfcc_data_o[113]));
 TIELOx1_ASAP7_75t_R _12890__115 (.L(mfcc_data_o[114]));
 TIELOx1_ASAP7_75t_R _12891__116 (.L(mfcc_data_o[115]));
 TIELOx1_ASAP7_75t_R _12892__117 (.L(mfcc_data_o[116]));
 TIELOx1_ASAP7_75t_R _12893__118 (.L(mfcc_data_o[117]));
 TIELOx1_ASAP7_75t_R _12894__119 (.L(mfcc_data_o[118]));
 TIELOx1_ASAP7_75t_R _12895__120 (.L(mfcc_data_o[119]));
 TIELOx1_ASAP7_75t_R _12896__121 (.L(mfcc_data_o[120]));
 TIELOx1_ASAP7_75t_R _12897__122 (.L(mfcc_data_o[121]));
 TIELOx1_ASAP7_75t_R _12898__123 (.L(mfcc_data_o[122]));
 TIELOx1_ASAP7_75t_R _12899__124 (.L(mfcc_data_o[123]));
 TIELOx1_ASAP7_75t_R _12900__125 (.L(mfcc_data_o[124]));
 TIELOx1_ASAP7_75t_R _12901__126 (.L(mfcc_data_o[125]));
 TIELOx1_ASAP7_75t_R _12902__127 (.L(mfcc_data_o[126]));
 TIELOx1_ASAP7_75t_R _12903__128 (.L(mfcc_data_o[127]));
 TIELOx1_ASAP7_75t_R _12904__129 (.L(mfcc_data_o[128]));
 TIELOx1_ASAP7_75t_R _12905__130 (.L(mfcc_data_o[129]));
 TIELOx1_ASAP7_75t_R _12906__131 (.L(mfcc_data_o[130]));
 TIELOx1_ASAP7_75t_R _12907__132 (.L(mfcc_data_o[131]));
 TIELOx1_ASAP7_75t_R _12908__133 (.L(mfcc_data_o[132]));
 TIELOx1_ASAP7_75t_R _12909__134 (.L(mfcc_data_o[133]));
 TIELOx1_ASAP7_75t_R _12910__135 (.L(mfcc_data_o[134]));
 TIELOx1_ASAP7_75t_R _12911__136 (.L(mfcc_data_o[135]));
 TIELOx1_ASAP7_75t_R _12912__137 (.L(mfcc_data_o[136]));
 TIELOx1_ASAP7_75t_R _12913__138 (.L(mfcc_data_o[137]));
 TIELOx1_ASAP7_75t_R _12914__139 (.L(mfcc_data_o[138]));
 TIELOx1_ASAP7_75t_R _12915__140 (.L(mfcc_data_o[139]));
 TIELOx1_ASAP7_75t_R _12916__141 (.L(mfcc_data_o[140]));
 TIELOx1_ASAP7_75t_R _12917__142 (.L(mfcc_data_o[141]));
 TIELOx1_ASAP7_75t_R _12918__143 (.L(mfcc_data_o[142]));
 TIELOx1_ASAP7_75t_R _12919__144 (.L(mfcc_data_o[143]));
 TIELOx1_ASAP7_75t_R _12920__145 (.L(mfcc_data_o[144]));
 TIELOx1_ASAP7_75t_R _12921__146 (.L(mfcc_data_o[145]));
 TIELOx1_ASAP7_75t_R _12922__147 (.L(mfcc_data_o[146]));
 TIELOx1_ASAP7_75t_R _12923__148 (.L(mfcc_data_o[147]));
 TIELOx1_ASAP7_75t_R _12924__149 (.L(mfcc_data_o[148]));
 TIELOx1_ASAP7_75t_R _12925__150 (.L(mfcc_data_o[149]));
 TIELOx1_ASAP7_75t_R _12926__151 (.L(mfcc_data_o[150]));
 TIELOx1_ASAP7_75t_R _12927__152 (.L(mfcc_data_o[151]));
 TIELOx1_ASAP7_75t_R _12928__153 (.L(mfcc_data_o[152]));
 TIELOx1_ASAP7_75t_R _12929__154 (.L(mfcc_data_o[153]));
 TIELOx1_ASAP7_75t_R _12930__155 (.L(mfcc_data_o[154]));
 TIELOx1_ASAP7_75t_R _12931__156 (.L(mfcc_data_o[155]));
 TIELOx1_ASAP7_75t_R _12932__157 (.L(mfcc_data_o[156]));
 TIELOx1_ASAP7_75t_R _12933__158 (.L(mfcc_data_o[157]));
 TIELOx1_ASAP7_75t_R _12934__159 (.L(mfcc_data_o[158]));
 TIELOx1_ASAP7_75t_R _12935__160 (.L(mfcc_data_o[159]));
 TIELOx1_ASAP7_75t_R _12936__161 (.L(mfcc_data_o[160]));
 TIELOx1_ASAP7_75t_R _12937__162 (.L(mfcc_data_o[161]));
 TIELOx1_ASAP7_75t_R _12938__163 (.L(mfcc_data_o[162]));
 TIELOx1_ASAP7_75t_R _12939__164 (.L(mfcc_data_o[163]));
 TIELOx1_ASAP7_75t_R _12940__165 (.L(mfcc_data_o[164]));
 TIELOx1_ASAP7_75t_R _12941__166 (.L(mfcc_data_o[165]));
 TIELOx1_ASAP7_75t_R _12942__167 (.L(mfcc_data_o[166]));
 TIELOx1_ASAP7_75t_R _12943__168 (.L(mfcc_data_o[167]));
 TIELOx1_ASAP7_75t_R _12944__169 (.L(mfcc_data_o[168]));
 TIELOx1_ASAP7_75t_R _12945__170 (.L(mfcc_data_o[169]));
 TIELOx1_ASAP7_75t_R _12946__171 (.L(mfcc_data_o[170]));
 TIELOx1_ASAP7_75t_R _12947__172 (.L(mfcc_data_o[171]));
 TIELOx1_ASAP7_75t_R _12948__173 (.L(mfcc_data_o[172]));
 TIELOx1_ASAP7_75t_R _12949__174 (.L(mfcc_data_o[173]));
 TIELOx1_ASAP7_75t_R _12950__175 (.L(mfcc_data_o[174]));
 TIELOx1_ASAP7_75t_R _12951__176 (.L(mfcc_data_o[175]));
 TIELOx1_ASAP7_75t_R _12952__177 (.L(mfcc_data_o[176]));
 TIELOx1_ASAP7_75t_R _12953__178 (.L(mfcc_data_o[177]));
 TIELOx1_ASAP7_75t_R _12954__179 (.L(mfcc_data_o[178]));
 TIELOx1_ASAP7_75t_R _12955__180 (.L(mfcc_data_o[179]));
 TIELOx1_ASAP7_75t_R _12956__181 (.L(mfcc_data_o[180]));
 TIELOx1_ASAP7_75t_R _12957__182 (.L(mfcc_data_o[181]));
 TIELOx1_ASAP7_75t_R _12958__183 (.L(mfcc_data_o[182]));
 TIELOx1_ASAP7_75t_R _12959__184 (.L(mfcc_data_o[183]));
 TIELOx1_ASAP7_75t_R _12960__185 (.L(mfcc_data_o[184]));
 TIELOx1_ASAP7_75t_R _12961__186 (.L(mfcc_data_o[185]));
 TIELOx1_ASAP7_75t_R _12962__187 (.L(mfcc_data_o[186]));
 TIELOx1_ASAP7_75t_R _12963__188 (.L(mfcc_data_o[187]));
 TIELOx1_ASAP7_75t_R _12964__189 (.L(mfcc_data_o[188]));
 TIELOx1_ASAP7_75t_R _12965__190 (.L(mfcc_data_o[189]));
 TIELOx1_ASAP7_75t_R _12966__191 (.L(mfcc_data_o[190]));
 TIELOx1_ASAP7_75t_R _12967__192 (.L(mfcc_data_o[191]));
 TIELOx1_ASAP7_75t_R _12968__193 (.L(mfcc_data_o[192]));
 TIELOx1_ASAP7_75t_R _12969__194 (.L(mfcc_data_o[193]));
 TIELOx1_ASAP7_75t_R _12970__195 (.L(mfcc_data_o[194]));
 TIELOx1_ASAP7_75t_R _12971__196 (.L(mfcc_data_o[195]));
 TIELOx1_ASAP7_75t_R _12972__197 (.L(mfcc_data_o[196]));
 TIELOx1_ASAP7_75t_R _12973__198 (.L(mfcc_data_o[197]));
 TIELOx1_ASAP7_75t_R _12974__199 (.L(mfcc_data_o[198]));
 TIELOx1_ASAP7_75t_R _12975__200 (.L(mfcc_data_o[199]));
 TIELOx1_ASAP7_75t_R _12976__201 (.L(mfcc_data_o[200]));
 TIELOx1_ASAP7_75t_R _12977__202 (.L(mfcc_data_o[201]));
 TIELOx1_ASAP7_75t_R _12978__203 (.L(mfcc_data_o[202]));
 TIELOx1_ASAP7_75t_R _12979__204 (.L(mfcc_data_o[203]));
 TIELOx1_ASAP7_75t_R _12980__205 (.L(mfcc_data_o[204]));
 TIELOx1_ASAP7_75t_R _12981__206 (.L(mfcc_data_o[205]));
 TIELOx1_ASAP7_75t_R _12982__207 (.L(mfcc_data_o[206]));
 TIELOx1_ASAP7_75t_R _12983__208 (.L(mfcc_data_o[207]));
 BUFx3_ASAP7_75t_R place3056 (.A(_06249_),
    .Y(net3056));
 BUFx3_ASAP7_75t_R place3057 (.A(_06243_),
    .Y(net3057));
 BUFx3_ASAP7_75t_R place3061 (.A(net5924),
    .Y(net3061));
 BUFx3_ASAP7_75t_R place3060 (.A(net5621),
    .Y(net3060));
 BUFx6f_ASAP7_75t_R place3062 (.A(_05143_),
    .Y(net3062));
 BUFx3_ASAP7_75t_R place3089 (.A(_06202_),
    .Y(net3089));
 BUFx3_ASAP7_75t_R place3066 (.A(_03911_),
    .Y(net3066));
 BUFx3_ASAP7_75t_R place3067 (.A(_03902_),
    .Y(net3067));
 BUFx3_ASAP7_75t_R place3068 (.A(_03896_),
    .Y(net3068));
 BUFx3_ASAP7_75t_R place3069 (.A(_02211_),
    .Y(net3069));
 BUFx3_ASAP7_75t_R place3070 (.A(_02195_),
    .Y(net3070));
 BUFx3_ASAP7_75t_R place3071 (.A(_02188_),
    .Y(net3071));
 BUFx3_ASAP7_75t_R place3072 (.A(_02175_),
    .Y(net3072));
 BUFx3_ASAP7_75t_R place3073 (.A(_02169_),
    .Y(net3073));
 BUFx3_ASAP7_75t_R place3074 (.A(_06261_),
    .Y(net3074));
 BUFx3_ASAP7_75t_R place3075 (.A(_06224_),
    .Y(net3075));
 BUFx3_ASAP7_75t_R place3076 (.A(_05142_),
    .Y(net3076));
 BUFx3_ASAP7_75t_R place3077 (.A(_05125_),
    .Y(net3077));
 BUFx3_ASAP7_75t_R place3078 (.A(_05097_),
    .Y(net3078));
 BUFx3_ASAP7_75t_R place3079 (.A(_03910_),
    .Y(net3079));
 BUFx3_ASAP7_75t_R place3080 (.A(_02192_),
    .Y(net3080));
 BUFx3_ASAP7_75t_R place3081 (.A(_02178_),
    .Y(net3081));
 BUFx3_ASAP7_75t_R place3082 (.A(_02174_),
    .Y(net3082));
 BUFx3_ASAP7_75t_R place3083 (.A(net5449),
    .Y(net3083));
 BUFx3_ASAP7_75t_R place3084 (.A(_02157_),
    .Y(net3084));
 BUFx3_ASAP7_75t_R place3085 (.A(_06236_),
    .Y(net3085));
 BUFx3_ASAP7_75t_R place3086 (.A(_06223_),
    .Y(net3086));
 BUFx3_ASAP7_75t_R place3087 (.A(_06214_),
    .Y(net3087));
 BUFx3_ASAP7_75t_R place3088 (.A(_06202_),
    .Y(net3088));
 BUFx3_ASAP7_75t_R place3090 (.A(_05130_),
    .Y(net3090));
 BUFx3_ASAP7_75t_R place3091 (.A(_05124_),
    .Y(net3091));
 BUFx3_ASAP7_75t_R place3092 (.A(_05111_),
    .Y(net3092));
 BUFx3_ASAP7_75t_R place3093 (.A(_05096_),
    .Y(net3093));
 BUFx3_ASAP7_75t_R place3094 (.A(_05085_),
    .Y(net3094));
 BUFx3_ASAP7_75t_R place3096 (.A(_02183_),
    .Y(net3096));
 BUFx3_ASAP7_75t_R place3097 (.A(_06242_),
    .Y(net3097));
 BUFx3_ASAP7_75t_R place3098 (.A(_06208_),
    .Y(net3098));
 BUFx3_ASAP7_75t_R place3099 (.A(_06197_),
    .Y(net3099));
 BUFx3_ASAP7_75t_R place3100 (.A(_05122_),
    .Y(net3100));
 BUFx3_ASAP7_75t_R place3102 (.A(_05087_),
    .Y(net3102));
 BUFx3_ASAP7_75t_R place3103 (.A(_03899_),
    .Y(net3103));
 BUFx3_ASAP7_75t_R place3104 (.A(_03893_),
    .Y(net3104));
 BUFx3_ASAP7_75t_R place3105 (.A(_03876_),
    .Y(net3105));
 BUFx3_ASAP7_75t_R place3106 (.A(_03871_),
    .Y(net3106));
 BUFx3_ASAP7_75t_R place3107 (.A(_02186_),
    .Y(net3107));
 BUFx3_ASAP7_75t_R place3108 (.A(_06227_),
    .Y(net3108));
 BUFx3_ASAP7_75t_R place3109 (.A(_06221_),
    .Y(net3109));
 BUFx3_ASAP7_75t_R place3110 (.A(_06207_),
    .Y(net3110));
 BUFx3_ASAP7_75t_R place3111 (.A(_06201_),
    .Y(net3111));
 BUFx3_ASAP7_75t_R place3112 (.A(net5663),
    .Y(net3112));
 BUFx3_ASAP7_75t_R place3113 (.A(net5627),
    .Y(net3113));
 BUFx3_ASAP7_75t_R place3114 (.A(_03875_),
    .Y(net3114));
 BUFx3_ASAP7_75t_R place3115 (.A(_03852_),
    .Y(net3115));
 BUFx3_ASAP7_75t_R place3116 (.A(_03835_),
    .Y(net3116));
 BUFx3_ASAP7_75t_R place3117 (.A(_02182_),
    .Y(net3117));
 BUFx3_ASAP7_75t_R place3119 (.A(_06210_),
    .Y(net3119));
 BUFx3_ASAP7_75t_R place3120 (.A(_06209_),
    .Y(net3120));
 BUFx3_ASAP7_75t_R place3121 (.A(_06204_),
    .Y(net3121));
 BUFx3_ASAP7_75t_R place3122 (.A(_06200_),
    .Y(net3122));
 BUFx3_ASAP7_75t_R place3123 (.A(_06194_),
    .Y(net3123));
 BUFx3_ASAP7_75t_R place3124 (.A(_05058_),
    .Y(net3124));
 BUFx3_ASAP7_75t_R place3125 (.A(_03834_),
    .Y(net3125));
 BUFx3_ASAP7_75t_R place3127 (.A(_02171_),
    .Y(net3127));
 BUFx3_ASAP7_75t_R place3128 (.A(_02134_),
    .Y(net3128));
 BUFx3_ASAP7_75t_R place3129 (.A(_02125_),
    .Y(net3129));
 BUFx6f_ASAP7_75t_R place3156 (.A(net3155),
    .Y(net3156));
 BUFx3_ASAP7_75t_R place3155 (.A(_03823_),
    .Y(net3155));
 BUFx3_ASAP7_75t_R place3132 (.A(_06192_),
    .Y(net3132));
 BUFx3_ASAP7_75t_R place3133 (.A(_06188_),
    .Y(net3133));
 BUFx3_ASAP7_75t_R place3142 (.A(net3141),
    .Y(net3142));
 BUFx3_ASAP7_75t_R place3134 (.A(_06183_),
    .Y(net3134));
 BUFx3_ASAP7_75t_R place3135 (.A(_05082_),
    .Y(net3135));
 BUFx3_ASAP7_75t_R place3136 (.A(_05076_),
    .Y(net3136));
 BUFx3_ASAP7_75t_R place3137 (.A(_05068_),
    .Y(net3137));
 BUFx3_ASAP7_75t_R place3138 (.A(_05055_),
    .Y(net3138));
 BUFx3_ASAP7_75t_R place3139 (.A(_05051_),
    .Y(net3139));
 BUFx3_ASAP7_75t_R place3140 (.A(net5972),
    .Y(net3140));
 BUFx3_ASAP7_75t_R place3141 (.A(_03858_),
    .Y(net3141));
 BUFx3_ASAP7_75t_R place3147 (.A(net3146),
    .Y(net3147));
 BUFx3_ASAP7_75t_R place3146 (.A(_06163_),
    .Y(net3146));
 BUFx3_ASAP7_75t_R place3143 (.A(_02140_),
    .Y(net3143));
 BUFx3_ASAP7_75t_R place3144 (.A(_02133_),
    .Y(net3144));
 BUFx3_ASAP7_75t_R place3145 (.A(_06186_),
    .Y(net3145));
 BUFx3_ASAP7_75t_R place3150 (.A(net3149),
    .Y(net3150));
 BUFx3_ASAP7_75t_R place3148 (.A(_06155_),
    .Y(net3148));
 BUFx6f_ASAP7_75t_R place3149 (.A(_05104_),
    .Y(net3149));
 BUFx3_ASAP7_75t_R place3151 (.A(_05081_),
    .Y(net3151));
 BUFx3_ASAP7_75t_R place3152 (.A(_05054_),
    .Y(net3152));
 BUFx3_ASAP7_75t_R place3153 (.A(_03843_),
    .Y(net3153));
 BUFx6f_ASAP7_75t_R place3154 (.A(_03826_),
    .Y(net3154));
 BUFx3_ASAP7_75t_R place3157 (.A(_02114_),
    .Y(net3157));
 BUFx3_ASAP7_75t_R place3158 (.A(_06195_),
    .Y(net3158));
 BUFx3_ASAP7_75t_R place3159 (.A(_06182_),
    .Y(net3159));
 BUFx3_ASAP7_75t_R place3162 (.A(_06154_),
    .Y(net3162));
 BUFx3_ASAP7_75t_R place3163 (.A(_05092_),
    .Y(net3163));
 BUFx3_ASAP7_75t_R place3164 (.A(_05061_),
    .Y(net3164));
 BUFx3_ASAP7_75t_R place3165 (.A(_03866_),
    .Y(net3165));
 BUFx3_ASAP7_75t_R place3166 (.A(net5681),
    .Y(net3166));
 BUFx3_ASAP7_75t_R place3168 (.A(_02147_),
    .Y(net3168));
 BUFx3_ASAP7_75t_R place3169 (.A(_02144_),
    .Y(net3169));
 BUFx3_ASAP7_75t_R place3170 (.A(_02131_),
    .Y(net3170));
 BUFx3_ASAP7_75t_R place3171 (.A(_02123_),
    .Y(net3171));
 BUFx3_ASAP7_75t_R place3172 (.A(_02101_),
    .Y(net3172));
 BUFx3_ASAP7_75t_R place3173 (.A(_02077_),
    .Y(net3173));
 BUFx3_ASAP7_75t_R place3174 (.A(_06159_),
    .Y(net3174));
 BUFx3_ASAP7_75t_R place3175 (.A(_06158_),
    .Y(net3175));
 BUFx3_ASAP7_75t_R place3176 (.A(net5936),
    .Y(net3176));
 BUFx3_ASAP7_75t_R place3178 (.A(_05064_),
    .Y(net3178));
 BUFx3_ASAP7_75t_R place3179 (.A(_03868_),
    .Y(net3179));
 BUFx3_ASAP7_75t_R place3180 (.A(_03862_),
    .Y(net3180));
 BUFx3_ASAP7_75t_R place3181 (.A(net5396),
    .Y(net3181));
 BUFx3_ASAP7_75t_R place3182 (.A(_02121_),
    .Y(net3182));
 BUFx3_ASAP7_75t_R place3183 (.A(_02111_),
    .Y(net3183));
 BUFx3_ASAP7_75t_R place3184 (.A(_02086_),
    .Y(net3184));
 BUFx3_ASAP7_75t_R place3190 (.A(_03800_),
    .Y(net3190));
 BUFx6f_ASAP7_75t_R place3185 (.A(_06130_),
    .Y(net3185));
 BUFx3_ASAP7_75t_R place3186 (.A(_05079_),
    .Y(net3186));
 BUFx3_ASAP7_75t_R place3187 (.A(_05041_),
    .Y(net3187));
 BUFx3_ASAP7_75t_R place3188 (.A(_05008_),
    .Y(net3188));
 BUFx3_ASAP7_75t_R place3189 (.A(_03822_),
    .Y(net3189));
 BUFx3_ASAP7_75t_R place3191 (.A(_03789_),
    .Y(net3191));
 BUFx3_ASAP7_75t_R place3192 (.A(_02129_),
    .Y(net3192));
 BUFx3_ASAP7_75t_R place3193 (.A(_02108_),
    .Y(net3193));
 BUFx3_ASAP7_75t_R place3194 (.A(_06135_),
    .Y(net3194));
 BUFx3_ASAP7_75t_R place3198 (.A(_05065_),
    .Y(net3198));
 BUFx3_ASAP7_75t_R place3199 (.A(_05046_),
    .Y(net3199));
 BUFx3_ASAP7_75t_R place3211 (.A(_06141_),
    .Y(net3211));
 BUFx3_ASAP7_75t_R place3200 (.A(_05023_),
    .Y(net3200));
 BUFx3_ASAP7_75t_R place3201 (.A(_05007_),
    .Y(net3201));
 BUFx3_ASAP7_75t_R place3202 (.A(_03819_),
    .Y(net3202));
 BUFx3_ASAP7_75t_R place3203 (.A(_03815_),
    .Y(net3203));
 BUFx3_ASAP7_75t_R place3204 (.A(_03799_),
    .Y(net3204));
 BUFx3_ASAP7_75t_R place3205 (.A(_03786_),
    .Y(net3205));
 BUFx3_ASAP7_75t_R place3206 (.A(_02097_),
    .Y(net3206));
 BUFx3_ASAP7_75t_R place3208 (.A(_06160_),
    .Y(net3208));
 BUFx6f_ASAP7_75t_R place3207 (.A(_06160_),
    .Y(net3207));
 BUFx3_ASAP7_75t_R place3209 (.A(_06150_),
    .Y(net3209));
 BUFx3_ASAP7_75t_R place3210 (.A(_06145_),
    .Y(net3210));
 BUFx3_ASAP7_75t_R place3213 (.A(_06108_),
    .Y(net3213));
 BUFx3_ASAP7_75t_R place3214 (.A(_05037_),
    .Y(net3214));
 BUFx3_ASAP7_75t_R place3215 (.A(_05027_),
    .Y(net3215));
 BUFx3_ASAP7_75t_R place3216 (.A(_05026_),
    .Y(net3216));
 BUFx3_ASAP7_75t_R place3217 (.A(_03805_),
    .Y(net3217));
 BUFx3_ASAP7_75t_R place3218 (.A(_03796_),
    .Y(net3218));
 BUFx3_ASAP7_75t_R place3219 (.A(_03787_),
    .Y(net3219));
 BUFx3_ASAP7_75t_R place3220 (.A(_02096_),
    .Y(net3220));
 BUFx3_ASAP7_75t_R place3221 (.A(_02094_),
    .Y(net3221));
 BUFx6f_ASAP7_75t_R place3222 (.A(_02071_),
    .Y(net3222));
 BUFx3_ASAP7_75t_R place3225 (.A(_06127_),
    .Y(net3225));
 BUFx3_ASAP7_75t_R place3223 (.A(net5443),
    .Y(net3223));
 BUFx3_ASAP7_75t_R place3224 (.A(_06144_),
    .Y(net3224));
 BUFx3_ASAP7_75t_R place3226 (.A(_06117_),
    .Y(net3226));
 BUFx3_ASAP7_75t_R place3227 (.A(_06107_),
    .Y(net3227));
 BUFx3_ASAP7_75t_R place3228 (.A(_05030_),
    .Y(net3228));
 BUFx3_ASAP7_75t_R place3230 (.A(_05005_),
    .Y(net3230));
 BUFx3_ASAP7_75t_R place3232 (.A(_03795_),
    .Y(net3232));
 BUFx3_ASAP7_75t_R place3233 (.A(net5980),
    .Y(net3233));
 BUFx3_ASAP7_75t_R place3234 (.A(net5669),
    .Y(net3234));
 BUFx3_ASAP7_75t_R place3235 (.A(_02092_),
    .Y(net3235));
 BUFx3_ASAP7_75t_R place3236 (.A(_02081_),
    .Y(net3236));
 BUFx3_ASAP7_75t_R place3237 (.A(_06143_),
    .Y(net3237));
 BUFx3_ASAP7_75t_R place3239 (.A(net5633),
    .Y(net3239));
 BUFx3_ASAP7_75t_R place3240 (.A(_05028_),
    .Y(net3240));
 BUFx3_ASAP7_75t_R place3241 (.A(_05001_),
    .Y(net3241));
 BUFx3_ASAP7_75t_R place3243 (.A(_03776_),
    .Y(net3243));
 BUFx3_ASAP7_75t_R place3245 (.A(_02075_),
    .Y(net3245));
 BUFx3_ASAP7_75t_R place3255 (.A(_05000_),
    .Y(net3255));
 BUFx3_ASAP7_75t_R place3248 (.A(_02069_),
    .Y(net3248));
 BUFx3_ASAP7_75t_R place3249 (.A(_02068_),
    .Y(net3249));
 BUFx3_ASAP7_75t_R place3250 (.A(_02038_),
    .Y(net3250));
 BUFx3_ASAP7_75t_R place3251 (.A(_06101_),
    .Y(net3251));
 BUFx3_ASAP7_75t_R place3252 (.A(_05019_),
    .Y(net3252));
 BUFx3_ASAP7_75t_R place3253 (.A(_05004_),
    .Y(net3253));
 BUFx3_ASAP7_75t_R place3254 (.A(_05003_),
    .Y(net3254));
 BUFx3_ASAP7_75t_R place3256 (.A(_04996_),
    .Y(net3256));
 BUFx3_ASAP7_75t_R place3257 (.A(_04988_),
    .Y(net3257));
 BUFx3_ASAP7_75t_R place3259 (.A(_04981_),
    .Y(net3259));
 BUFx3_ASAP7_75t_R place3260 (.A(_04974_),
    .Y(net3260));
 BUFx3_ASAP7_75t_R place3261 (.A(_04965_),
    .Y(net3261));
 BUFx3_ASAP7_75t_R place3262 (.A(net5998),
    .Y(net3262));
 BUFx3_ASAP7_75t_R place3263 (.A(_03767_),
    .Y(net3263));
 BUFx3_ASAP7_75t_R place3264 (.A(_03760_),
    .Y(net3264));
 BUFx3_ASAP7_75t_R place3266 (.A(_02090_),
    .Y(net3266));
 BUFx3_ASAP7_75t_R place3268 (.A(_06099_),
    .Y(net3268));
 BUFx6f_ASAP7_75t_R place3269 (.A(_06097_),
    .Y(net3269));
 BUFx3_ASAP7_75t_R place3270 (.A(_06088_),
    .Y(net3270));
 BUFx3_ASAP7_75t_R place3271 (.A(_04976_),
    .Y(net3271));
 BUFx3_ASAP7_75t_R place3272 (.A(_04964_),
    .Y(net3272));
 BUFx3_ASAP7_75t_R place3273 (.A(_04946_),
    .Y(net3273));
 BUFx3_ASAP7_75t_R place3274 (.A(_03759_),
    .Y(net3274));
 BUFx3_ASAP7_75t_R place3275 (.A(_03736_),
    .Y(net3275));
 BUFx3_ASAP7_75t_R place3281 (.A(_06118_),
    .Y(net3281));
 BUFx3_ASAP7_75t_R place3277 (.A(_02089_),
    .Y(net3277));
 BUFx3_ASAP7_75t_R place3278 (.A(_02059_),
    .Y(net3278));
 BUFx3_ASAP7_75t_R place3279 (.A(_02047_),
    .Y(net3279));
 BUFx3_ASAP7_75t_R place3280 (.A(_02028_),
    .Y(net3280));
 BUFx3_ASAP7_75t_R place3282 (.A(_06112_),
    .Y(net3282));
 BUFx3_ASAP7_75t_R place3283 (.A(_06104_),
    .Y(net3283));
 BUFx3_ASAP7_75t_R place3284 (.A(_06096_),
    .Y(net3284));
 BUFx3_ASAP7_75t_R place3285 (.A(net5625),
    .Y(net3285));
 BUFx3_ASAP7_75t_R place3286 (.A(_06058_),
    .Y(net3286));
 BUFx3_ASAP7_75t_R place3287 (.A(_04972_),
    .Y(net3287));
 BUFx3_ASAP7_75t_R place3288 (.A(_04963_),
    .Y(net3288));
 BUFx3_ASAP7_75t_R place3294 (.A(_03741_),
    .Y(net3294));
 BUFx3_ASAP7_75t_R place3289 (.A(_03771_),
    .Y(net3289));
 BUFx3_ASAP7_75t_R place3290 (.A(_03763_),
    .Y(net3290));
 BUFx3_ASAP7_75t_R place3291 (.A(_03758_),
    .Y(net3291));
 BUFx3_ASAP7_75t_R place3292 (.A(net5703),
    .Y(net3292));
 BUFx3_ASAP7_75t_R place3293 (.A(_03741_),
    .Y(net3293));
 BUFx3_ASAP7_75t_R place3322 (.A(_02004_),
    .Y(net3322));
 BUFx3_ASAP7_75t_R place3295 (.A(_02066_),
    .Y(net3295));
 BUFx3_ASAP7_75t_R place3296 (.A(net5765),
    .Y(net3296));
 BUFx3_ASAP7_75t_R place3297 (.A(_02046_),
    .Y(net3297));
 BUFx3_ASAP7_75t_R place3298 (.A(net5442),
    .Y(net3298));
 BUFx3_ASAP7_75t_R place3299 (.A(_02027_),
    .Y(net3299));
 BUFx3_ASAP7_75t_R place3300 (.A(_02022_),
    .Y(net3300));
 BUFx3_ASAP7_75t_R place3301 (.A(_02007_),
    .Y(net3301));
 BUFx3_ASAP7_75t_R place3302 (.A(_06092_),
    .Y(net3302));
 BUFx3_ASAP7_75t_R place3303 (.A(_06077_),
    .Y(net3303));
 BUFx3_ASAP7_75t_R place3304 (.A(_04983_),
    .Y(net3304));
 BUFx3_ASAP7_75t_R place3305 (.A(_04977_),
    .Y(net3305));
 BUFx3_ASAP7_75t_R place3306 (.A(_04971_),
    .Y(net3306));
 BUFx3_ASAP7_75t_R place3307 (.A(_04962_),
    .Y(net3307));
 BUFx3_ASAP7_75t_R place3308 (.A(_04956_),
    .Y(net3308));
 BUFx3_ASAP7_75t_R place3309 (.A(_04952_),
    .Y(net3309));
 BUFx3_ASAP7_75t_R place3310 (.A(_04941_),
    .Y(net3310));
 BUFx3_ASAP7_75t_R place3311 (.A(_04925_),
    .Y(net3311));
 BUFx3_ASAP7_75t_R place3318 (.A(net3317),
    .Y(net3318));
 BUFx3_ASAP7_75t_R place3312 (.A(_03756_),
    .Y(net3312));
 BUFx3_ASAP7_75t_R place3313 (.A(net5694),
    .Y(net3313));
 BUFx3_ASAP7_75t_R place3314 (.A(_03745_),
    .Y(net3314));
 BUFx3_ASAP7_75t_R place3315 (.A(_03729_),
    .Y(net3315));
 BUFx3_ASAP7_75t_R place3316 (.A(_02043_),
    .Y(net3316));
 BUFx6f_ASAP7_75t_R place3317 (.A(_02042_),
    .Y(net3317));
 BUFx3_ASAP7_75t_R place3319 (.A(net5387),
    .Y(net3319));
 BUFx3_ASAP7_75t_R place3320 (.A(_02030_),
    .Y(net3320));
 BUFx3_ASAP7_75t_R place3321 (.A(_02004_),
    .Y(net3321));
 BUFx3_ASAP7_75t_R place3323 (.A(_06091_),
    .Y(net3323));
 BUFx3_ASAP7_75t_R place3324 (.A(_04970_),
    .Y(net3324));
 BUFx3_ASAP7_75t_R place3326 (.A(_04948_),
    .Y(net3326));
 BUFx3_ASAP7_75t_R place3327 (.A(_04931_),
    .Y(net3327));
 BUFx3_ASAP7_75t_R place3328 (.A(_04924_),
    .Y(net3328));
 BUFx3_ASAP7_75t_R place3329 (.A(_03808_),
    .Y(net3329));
 BUFx3_ASAP7_75t_R place3330 (.A(_03765_),
    .Y(net3330));
 BUFx3_ASAP7_75t_R place3332 (.A(_03728_),
    .Y(net3332));
 BUFx6f_ASAP7_75t_R place3334 (.A(_03719_),
    .Y(net3334));
 BUFx3_ASAP7_75t_R place3343 (.A(_04938_),
    .Y(net3343));
 BUFx3_ASAP7_75t_R place3336 (.A(_02044_),
    .Y(net3336));
 BUFx3_ASAP7_75t_R place3337 (.A(_02005_),
    .Y(net3337));
 BUFx3_ASAP7_75t_R place3338 (.A(_01991_),
    .Y(net3338));
 BUFx3_ASAP7_75t_R place3339 (.A(_06063_),
    .Y(net3339));
 BUFx3_ASAP7_75t_R place3340 (.A(_06045_),
    .Y(net3340));
 BUFx3_ASAP7_75t_R place3341 (.A(_06030_),
    .Y(net3341));
 BUFx3_ASAP7_75t_R place3342 (.A(_04938_),
    .Y(net3342));
 BUFx3_ASAP7_75t_R place3344 (.A(_04909_),
    .Y(net3344));
 BUFx3_ASAP7_75t_R place3453 (.A(_05981_),
    .Y(net3453));
 BUFx3_ASAP7_75t_R place3345 (.A(_03742_),
    .Y(net3345));
 BUFx3_ASAP7_75t_R place3349 (.A(net3348),
    .Y(net3349));
 BUFx3_ASAP7_75t_R place3346 (.A(net5682),
    .Y(net3346));
 BUFx3_ASAP7_75t_R place3347 (.A(_03718_),
    .Y(net3347));
 BUFx6f_ASAP7_75t_R place3348 (.A(_03706_),
    .Y(net3348));
 BUFx3_ASAP7_75t_R place3448 (.A(net5424),
    .Y(net3448));
 BUFx3_ASAP7_75t_R place3378 (.A(_01963_),
    .Y(net3378));
 BUFx3_ASAP7_75t_R place3350 (.A(_02018_),
    .Y(net3350));
 BUFx3_ASAP7_75t_R place3351 (.A(_02015_),
    .Y(net3351));
 BUFx3_ASAP7_75t_R place3352 (.A(net5422),
    .Y(net3352));
 BUFx3_ASAP7_75t_R place3353 (.A(net5773),
    .Y(net3353));
 BUFx3_ASAP7_75t_R place3354 (.A(_01990_),
    .Y(net3354));
 BUFx3_ASAP7_75t_R place3355 (.A(_01979_),
    .Y(net3355));
 BUFx3_ASAP7_75t_R place3356 (.A(_06067_),
    .Y(net3356));
 BUFx3_ASAP7_75t_R place3357 (.A(net5624),
    .Y(net3357));
 BUFx3_ASAP7_75t_R place3358 (.A(_06044_),
    .Y(net3358));
 BUFx3_ASAP7_75t_R place3359 (.A(_06040_),
    .Y(net3359));
 BUFx3_ASAP7_75t_R place3360 (.A(_04958_),
    .Y(net3360));
 BUFx3_ASAP7_75t_R place3361 (.A(_03732_),
    .Y(net3361));
 BUFx3_ASAP7_75t_R place3362 (.A(_03731_),
    .Y(net3362));
 BUFx3_ASAP7_75t_R place3363 (.A(net5700),
    .Y(net3363));
 BUFx3_ASAP7_75t_R place3364 (.A(_03714_),
    .Y(net3364));
 BUFx6f_ASAP7_75t_R place3365 (.A(_03686_),
    .Y(net3365));
 BUFx3_ASAP7_75t_R place3366 (.A(_02009_),
    .Y(net3366));
 BUFx3_ASAP7_75t_R place3367 (.A(_02002_),
    .Y(net3367));
 BUFx3_ASAP7_75t_R place3368 (.A(_06089_),
    .Y(net3368));
 BUFx3_ASAP7_75t_R place3369 (.A(_06064_),
    .Y(net3369));
 BUFx3_ASAP7_75t_R place3370 (.A(_04957_),
    .Y(net3370));
 BUFx3_ASAP7_75t_R place3371 (.A(_04927_),
    .Y(net3371));
 BUFx3_ASAP7_75t_R place3372 (.A(_04921_),
    .Y(net3372));
 BUFx3_ASAP7_75t_R place3373 (.A(_04912_),
    .Y(net3373));
 BUFx3_ASAP7_75t_R place3374 (.A(_03725_),
    .Y(net3374));
 BUFx3_ASAP7_75t_R place3375 (.A(_01988_),
    .Y(net3375));
 BUFx3_ASAP7_75t_R place3376 (.A(_01977_),
    .Y(net3376));
 BUFx3_ASAP7_75t_R place3377 (.A(_01963_),
    .Y(net3377));
 BUFx3_ASAP7_75t_R place3430 (.A(_01933_),
    .Y(net3430));
 BUFx3_ASAP7_75t_R place3379 (.A(net5600),
    .Y(net3379));
 BUFx3_ASAP7_75t_R place3380 (.A(_06050_),
    .Y(net3380));
 BUFx3_ASAP7_75t_R place3425 (.A(net3424),
    .Y(net3425));
 BUFx3_ASAP7_75t_R place3381 (.A(_04934_),
    .Y(net3381));
 BUFx3_ASAP7_75t_R place3382 (.A(_04917_),
    .Y(net3382));
 BUFx6f_ASAP7_75t_R place3383 (.A(_04911_),
    .Y(net3383));
 BUFx3_ASAP7_75t_R place3384 (.A(_04903_),
    .Y(net3384));
 BUFx3_ASAP7_75t_R place3385 (.A(_04891_),
    .Y(net3385));
 BUFx3_ASAP7_75t_R place3386 (.A(_04888_),
    .Y(net3386));
 BUFx3_ASAP7_75t_R place3387 (.A(_03721_),
    .Y(net3387));
 BUFx3_ASAP7_75t_R place3388 (.A(_03697_),
    .Y(net3388));
 BUFx3_ASAP7_75t_R place3389 (.A(_03680_),
    .Y(net3389));
 BUFx3_ASAP7_75t_R place3390 (.A(_03671_),
    .Y(net3390));
 BUFx3_ASAP7_75t_R place3391 (.A(_01987_),
    .Y(net3391));
 BUFx6f_ASAP7_75t_R place3392 (.A(_01962_),
    .Y(net3392));
 BUFx3_ASAP7_75t_R place3393 (.A(_06037_),
    .Y(net3393));
 BUFx3_ASAP7_75t_R place3394 (.A(_03696_),
    .Y(net3394));
 BUFx3_ASAP7_75t_R place3395 (.A(_03690_),
    .Y(net3395));
 BUFx3_ASAP7_75t_R place3396 (.A(net5988),
    .Y(net3396));
 BUFx3_ASAP7_75t_R place3397 (.A(_03679_),
    .Y(net3397));
 BUFx3_ASAP7_75t_R place3398 (.A(_03670_),
    .Y(net3398));
 BUFx3_ASAP7_75t_R place3400 (.A(net5996),
    .Y(net3400));
 BUFx3_ASAP7_75t_R place3399 (.A(_03651_),
    .Y(net3399));
 BUFx3_ASAP7_75t_R place3422 (.A(_04866_),
    .Y(net3422));
 BUFx3_ASAP7_75t_R place3401 (.A(_01986_),
    .Y(net3401));
 BUFx3_ASAP7_75t_R place3402 (.A(_01971_),
    .Y(net3402));
 BUFx3_ASAP7_75t_R place3403 (.A(_01961_),
    .Y(net3403));
 BUFx3_ASAP7_75t_R place3404 (.A(_01957_),
    .Y(net3404));
 BUFx3_ASAP7_75t_R place3405 (.A(net5423),
    .Y(net3405));
 BUFx3_ASAP7_75t_R place3408 (.A(_06017_),
    .Y(net3408));
 BUFx3_ASAP7_75t_R place3406 (.A(_06052_),
    .Y(net3406));
 BUFx3_ASAP7_75t_R place3407 (.A(_06024_),
    .Y(net3407));
 BUFx3_ASAP7_75t_R place3418 (.A(net3417),
    .Y(net3418));
 BUFx3_ASAP7_75t_R place3409 (.A(_06003_),
    .Y(net3409));
 BUFx3_ASAP7_75t_R place3413 (.A(_03660_),
    .Y(net3413));
 BUFx3_ASAP7_75t_R place3410 (.A(_04879_),
    .Y(net3410));
 BUFx3_ASAP7_75t_R place3411 (.A(_03700_),
    .Y(net3411));
 BUFx3_ASAP7_75t_R place3412 (.A(_03695_),
    .Y(net3412));
 BUFx3_ASAP7_75t_R place3414 (.A(_01966_),
    .Y(net3414));
 BUFx3_ASAP7_75t_R place3415 (.A(_01956_),
    .Y(net3415));
 BUFx3_ASAP7_75t_R place3416 (.A(_01948_),
    .Y(net3416));
 BUFx3_ASAP7_75t_R place3417 (.A(_01939_),
    .Y(net3417));
 BUFx3_ASAP7_75t_R place3419 (.A(_06021_),
    .Y(net3419));
 BUFx3_ASAP7_75t_R place3420 (.A(_06008_),
    .Y(net3420));
 BUFx3_ASAP7_75t_R place3421 (.A(_04913_),
    .Y(net3421));
 BUFx3_ASAP7_75t_R place3423 (.A(_03674_),
    .Y(net3423));
 BUFx3_ASAP7_75t_R place3424 (.A(_03668_),
    .Y(net3424));
 BUFx3_ASAP7_75t_R place3426 (.A(_03649_),
    .Y(net3426));
 BUFx3_ASAP7_75t_R place3427 (.A(_01959_),
    .Y(net3427));
 BUFx3_ASAP7_75t_R rebuffer5910 (.A(_04330_),
    .Y(net5910));
 BUFx3_ASAP7_75t_R place3429 (.A(_01935_),
    .Y(net3429));
 BUFx3_ASAP7_75t_R place3440 (.A(net3439),
    .Y(net3440));
 BUFx3_ASAP7_75t_R place3431 (.A(_06022_),
    .Y(net3431));
 BUFx3_ASAP7_75t_R place3432 (.A(_06009_),
    .Y(net3432));
 BUFx3_ASAP7_75t_R place3433 (.A(_05998_),
    .Y(net3433));
 BUFx3_ASAP7_75t_R place3434 (.A(_05983_),
    .Y(net3434));
 BUFx3_ASAP7_75t_R place3435 (.A(_04899_),
    .Y(net3435));
 BUFx3_ASAP7_75t_R place3436 (.A(_04896_),
    .Y(net3436));
 BUFx3_ASAP7_75t_R place3437 (.A(_04893_),
    .Y(net3437));
 BUFx3_ASAP7_75t_R place3438 (.A(_04885_),
    .Y(net3438));
 BUFx3_ASAP7_75t_R place3439 (.A(_04865_),
    .Y(net3439));
 BUFx3_ASAP7_75t_R place3441 (.A(_03673_),
    .Y(net3441));
 BUFx3_ASAP7_75t_R place3442 (.A(_03653_),
    .Y(net3442));
 BUFx3_ASAP7_75t_R place3443 (.A(_03645_),
    .Y(net3443));
 BUFx3_ASAP7_75t_R place3444 (.A(_01954_),
    .Y(net3444));
 BUFx3_ASAP7_75t_R place3445 (.A(_01953_),
    .Y(net3445));
 BUFx3_ASAP7_75t_R place3446 (.A(_01951_),
    .Y(net3446));
 BUFx3_ASAP7_75t_R place3447 (.A(net5424),
    .Y(net3447));
 BUFx3_ASAP7_75t_R place3449 (.A(_01927_),
    .Y(net3449));
 BUFx3_ASAP7_75t_R place3450 (.A(_01903_),
    .Y(net3450));
 BUFx3_ASAP7_75t_R place3451 (.A(_06001_),
    .Y(net3451));
 BUFx3_ASAP7_75t_R place3452 (.A(net5638),
    .Y(net3452));
 BUFx3_ASAP7_75t_R place3454 (.A(_04878_),
    .Y(net3454));
 BUFx3_ASAP7_75t_R place3455 (.A(_04869_),
    .Y(net3455));
 BUFx3_ASAP7_75t_R place3456 (.A(_03672_),
    .Y(net3456));
 BUFx3_ASAP7_75t_R place3457 (.A(net5982),
    .Y(net3457));
 BUFx3_ASAP7_75t_R place3458 (.A(_03647_),
    .Y(net3458));
 BUFx3_ASAP7_75t_R place3460 (.A(net5704),
    .Y(net3460));
 BUFx3_ASAP7_75t_R place3461 (.A(net5999),
    .Y(net3461));
 BUFx3_ASAP7_75t_R place3462 (.A(_03628_),
    .Y(net3462));
 BUFx3_ASAP7_75t_R place3533 (.A(_04829_),
    .Y(net3533));
 BUFx3_ASAP7_75t_R place3513 (.A(_05906_),
    .Y(net3513));
 BUFx3_ASAP7_75t_R place3506 (.A(_01876_),
    .Y(net3506));
 BUFx3_ASAP7_75t_R place3463 (.A(net5388),
    .Y(net3463));
 BUFx3_ASAP7_75t_R place3482 (.A(_03632_),
    .Y(net3482));
 BUFx3_ASAP7_75t_R place3469 (.A(_04870_),
    .Y(net3469));
 BUFx3_ASAP7_75t_R place3464 (.A(_01902_),
    .Y(net3464));
 BUFx3_ASAP7_75t_R place3465 (.A(_06023_),
    .Y(net3465));
 BUFx3_ASAP7_75t_R place3466 (.A(net5940),
    .Y(net3466));
 BUFx3_ASAP7_75t_R place3467 (.A(net5934),
    .Y(net3467));
 BUFx3_ASAP7_75t_R place3468 (.A(_05944_),
    .Y(net3468));
 BUFx3_ASAP7_75t_R place3470 (.A(_04854_),
    .Y(net3470));
 BUFx3_ASAP7_75t_R place3471 (.A(_03655_),
    .Y(net3471));
 BUFx3_ASAP7_75t_R place3472 (.A(_03654_),
    .Y(net3472));
 BUFx3_ASAP7_75t_R place3473 (.A(_03640_),
    .Y(net3473));
 BUFx3_ASAP7_75t_R place3474 (.A(_03634_),
    .Y(net3474));
 BUFx3_ASAP7_75t_R place3475 (.A(_01958_),
    .Y(net3475));
 BUFx3_ASAP7_75t_R place3476 (.A(_01886_),
    .Y(net3476));
 BUFx3_ASAP7_75t_R place3477 (.A(_06010_),
    .Y(net3477));
 BUFx3_ASAP7_75t_R place3478 (.A(_05964_),
    .Y(net3478));
 BUFx3_ASAP7_75t_R place3479 (.A(_05960_),
    .Y(net3479));
 BUFx3_ASAP7_75t_R place3480 (.A(_04863_),
    .Y(net3480));
 BUFx3_ASAP7_75t_R place3481 (.A(_03633_),
    .Y(net3481));
 BUFx6f_ASAP7_75t_R place3483 (.A(net5675),
    .Y(net3483));
 BUFx3_ASAP7_75t_R place3484 (.A(_01901_),
    .Y(net3484));
 BUFx3_ASAP7_75t_R place3485 (.A(_01885_),
    .Y(net3485));
 BUFx3_ASAP7_75t_R place3486 (.A(net5629),
    .Y(net3486));
 BUFx3_ASAP7_75t_R place3487 (.A(_05973_),
    .Y(net3487));
 BUFx3_ASAP7_75t_R place3488 (.A(_05940_),
    .Y(net3488));
 BUFx3_ASAP7_75t_R place3489 (.A(_04857_),
    .Y(net3489));
 BUFx3_ASAP7_75t_R place3490 (.A(_03625_),
    .Y(net3490));
 BUFx3_ASAP7_75t_R place3491 (.A(net5389),
    .Y(net3491));
 BUFx3_ASAP7_75t_R place3497 (.A(_04845_),
    .Y(net3497));
 BUFx3_ASAP7_75t_R place3492 (.A(_01884_),
    .Y(net3492));
 BUFx3_ASAP7_75t_R place3493 (.A(_05962_),
    .Y(net3493));
 BUFx3_ASAP7_75t_R place3494 (.A(_04872_),
    .Y(net3494));
 BUFx3_ASAP7_75t_R place3495 (.A(_04862_),
    .Y(net3495));
 BUFx3_ASAP7_75t_R place3496 (.A(_04851_),
    .Y(net3496));
 BUFx3_ASAP7_75t_R place3498 (.A(_04832_),
    .Y(net3498));
 BUFx3_ASAP7_75t_R place3499 (.A(_03635_),
    .Y(net3499));
 BUFx3_ASAP7_75t_R place3500 (.A(_03619_),
    .Y(net3500));
 BUFx3_ASAP7_75t_R place3501 (.A(net5997),
    .Y(net3501));
 BUFx3_ASAP7_75t_R place3502 (.A(_03609_),
    .Y(net3502));
 BUFx3_ASAP7_75t_R place3503 (.A(net5986),
    .Y(net3503));
 BUFx3_ASAP7_75t_R place3504 (.A(_03580_),
    .Y(net3504));
 BUFx3_ASAP7_75t_R place3505 (.A(_01898_),
    .Y(net3505));
 BUFx3_ASAP7_75t_R place3507 (.A(_05959_),
    .Y(net3507));
 BUFx3_ASAP7_75t_R place3508 (.A(_05952_),
    .Y(net3508));
 BUFx3_ASAP7_75t_R place3509 (.A(_05947_),
    .Y(net3509));
 BUFx3_ASAP7_75t_R place3510 (.A(_05938_),
    .Y(net3510));
 BUFx3_ASAP7_75t_R place3512 (.A(_05906_),
    .Y(net3512));
 BUFx6f_ASAP7_75t_R place3511 (.A(_05906_),
    .Y(net3511));
 BUFx6f_ASAP7_75t_R place3518 (.A(_01912_),
    .Y(net3518));
 BUFx3_ASAP7_75t_R place3514 (.A(_04871_),
    .Y(net3514));
 BUFx3_ASAP7_75t_R place3515 (.A(_04830_),
    .Y(net3515));
 BUFx3_ASAP7_75t_R place3516 (.A(_04810_),
    .Y(net3516));
 BUFx3_ASAP7_75t_R place3517 (.A(net5691),
    .Y(net3517));
 BUFx3_ASAP7_75t_R place3519 (.A(_01905_),
    .Y(net3519));
 BUFx3_ASAP7_75t_R place3520 (.A(_01900_),
    .Y(net3520));
 BUFx3_ASAP7_75t_R place3521 (.A(_01893_),
    .Y(net3521));
 BUFx3_ASAP7_75t_R place3522 (.A(_01882_),
    .Y(net3522));
 BUFx3_ASAP7_75t_R place3523 (.A(_05946_),
    .Y(net3523));
 BUFx3_ASAP7_75t_R place3524 (.A(_05945_),
    .Y(net3524));
 BUFx3_ASAP7_75t_R place3525 (.A(_05943_),
    .Y(net3525));
 BUFx3_ASAP7_75t_R place3526 (.A(_05937_),
    .Y(net3526));
 BUFx3_ASAP7_75t_R place3527 (.A(_05914_),
    .Y(net3527));
 BUFx3_ASAP7_75t_R place3528 (.A(_05905_),
    .Y(net3528));
 BUFx3_ASAP7_75t_R place3529 (.A(_04859_),
    .Y(net3529));
 BUFx3_ASAP7_75t_R place3530 (.A(_04858_),
    .Y(net3530));
 BUFx3_ASAP7_75t_R place3531 (.A(_04842_),
    .Y(net3531));
 BUFx3_ASAP7_75t_R place3532 (.A(_04831_),
    .Y(net3532));
 BUFx3_ASAP7_75t_R place3534 (.A(_04805_),
    .Y(net3534));
 BUFx3_ASAP7_75t_R place3536 (.A(net5667),
    .Y(net3536));
 BUFx3_ASAP7_75t_R place3537 (.A(_01897_),
    .Y(net3537));
 BUFx3_ASAP7_75t_R place3538 (.A(_01894_),
    .Y(net3538));
 BUFx3_ASAP7_75t_R place3539 (.A(_01892_),
    .Y(net3539));
 BUFx3_ASAP7_75t_R place3540 (.A(_01890_),
    .Y(net3540));
 BUFx6f_ASAP7_75t_R place3541 (.A(_01852_),
    .Y(net3541));
 BUFx3_ASAP7_75t_R place3542 (.A(_05936_),
    .Y(net3542));
 BUFx3_ASAP7_75t_R place3543 (.A(_05935_),
    .Y(net3543));
 BUFx3_ASAP7_75t_R place3544 (.A(_05927_),
    .Y(net3544));
 BUFx3_ASAP7_75t_R place3545 (.A(_05921_),
    .Y(net3545));
 BUFx3_ASAP7_75t_R place3546 (.A(_04840_),
    .Y(net3546));
 BUFx3_ASAP7_75t_R place3547 (.A(_04822_),
    .Y(net3547));
 BUFx3_ASAP7_75t_R place3549 (.A(_03575_),
    .Y(net3549));
 BUFx3_ASAP7_75t_R place3550 (.A(_03570_),
    .Y(net3550));
 BUFx3_ASAP7_75t_R place3551 (.A(_03558_),
    .Y(net3551));
 BUFx3_ASAP7_75t_R place3552 (.A(net5760),
    .Y(net3552));
 BUFx3_ASAP7_75t_R place3553 (.A(_01869_),
    .Y(net3553));
 BUFx3_ASAP7_75t_R place3560 (.A(_03593_),
    .Y(net3560));
 BUFx3_ASAP7_75t_R place3554 (.A(_05932_),
    .Y(net3554));
 BUFx3_ASAP7_75t_R place3555 (.A(_05920_),
    .Y(net3555));
 BUFx3_ASAP7_75t_R place3556 (.A(_05912_),
    .Y(net3556));
 BUFx3_ASAP7_75t_R place3557 (.A(_05903_),
    .Y(net3557));
 BUFx3_ASAP7_75t_R place3558 (.A(_04843_),
    .Y(net3558));
 BUFx3_ASAP7_75t_R place3559 (.A(_04795_),
    .Y(net3559));
 BUFx3_ASAP7_75t_R place3561 (.A(_03577_),
    .Y(net3561));
 BUFx3_ASAP7_75t_R place3562 (.A(net5705),
    .Y(net3562));
 BUFx3_ASAP7_75t_R place3563 (.A(_03569_),
    .Y(net3563));
 BUFx6f_ASAP7_75t_R rebuffer6001 (.A(_03435_),
    .Y(net6001));
 BUFx3_ASAP7_75t_R place3565 (.A(_01863_),
    .Y(net3565));
 BUFx3_ASAP7_75t_R place3566 (.A(_01826_),
    .Y(net3566));
 BUFx3_ASAP7_75t_R place3567 (.A(_05934_),
    .Y(net3567));
 BUFx3_ASAP7_75t_R place3568 (.A(_05929_),
    .Y(net3568));
 BUFx3_ASAP7_75t_R place3569 (.A(_05924_),
    .Y(net3569));
 BUFx3_ASAP7_75t_R place3570 (.A(net5935),
    .Y(net3570));
 BUFx3_ASAP7_75t_R place3571 (.A(_04802_),
    .Y(net3571));
 BUFx3_ASAP7_75t_R place3573 (.A(_04786_),
    .Y(net3573));
 BUFx3_ASAP7_75t_R place3574 (.A(_04777_),
    .Y(net3574));
 BUFx3_ASAP7_75t_R place3575 (.A(_03588_),
    .Y(net3575));
 BUFx3_ASAP7_75t_R place3577 (.A(net5973),
    .Y(net3577));
 BUFx3_ASAP7_75t_R place3578 (.A(_01879_),
    .Y(net3578));
 BUFx3_ASAP7_75t_R place3579 (.A(_01877_),
    .Y(net3579));
 BUFx3_ASAP7_75t_R place3580 (.A(_01872_),
    .Y(net3580));
 BUFx3_ASAP7_75t_R place3581 (.A(_01867_),
    .Y(net3581));
 BUFx3_ASAP7_75t_R place3582 (.A(_01862_),
    .Y(net3582));
 BUFx3_ASAP7_75t_R place3583 (.A(_01848_),
    .Y(net3583));
 BUFx3_ASAP7_75t_R place3584 (.A(_01842_),
    .Y(net3584));
 BUFx3_ASAP7_75t_R place3585 (.A(net5937),
    .Y(net3585));
 BUFx3_ASAP7_75t_R place3586 (.A(_05891_),
    .Y(net3586));
 BUFx3_ASAP7_75t_R place3587 (.A(_05886_),
    .Y(net3587));
 BUFx6f_ASAP7_75t_R place3588 (.A(_05881_),
    .Y(net3588));
 BUFx3_ASAP7_75t_R place3589 (.A(_04800_),
    .Y(net3589));
 BUFx3_ASAP7_75t_R place3591 (.A(_04774_),
    .Y(net3591));
 BUFx3_ASAP7_75t_R place3592 (.A(net5985),
    .Y(net3592));
 BUFx3_ASAP7_75t_R place3613 (.A(net3612),
    .Y(net3613));
 BUFx3_ASAP7_75t_R place3594 (.A(_03546_),
    .Y(net3594));
 BUFx3_ASAP7_75t_R place3595 (.A(_01851_),
    .Y(net3595));
 BUFx6f_ASAP7_75t_R place3596 (.A(_01837_),
    .Y(net3596));
 BUFx3_ASAP7_75t_R place3597 (.A(_01831_),
    .Y(net3597));
 BUFx3_ASAP7_75t_R place3603 (.A(_04798_),
    .Y(net3603));
 BUFx3_ASAP7_75t_R place3598 (.A(_04779_),
    .Y(net3598));
 BUFx3_ASAP7_75t_R place3599 (.A(_03552_),
    .Y(net3599));
 BUFx3_ASAP7_75t_R place3600 (.A(_03535_),
    .Y(net3600));
 BUFx3_ASAP7_75t_R place3601 (.A(_05867_),
    .Y(net3601));
 BUFx3_ASAP7_75t_R place3602 (.A(_05856_),
    .Y(net3602));
 BUFx3_ASAP7_75t_R place3604 (.A(_04783_),
    .Y(net3604));
 BUFx3_ASAP7_75t_R place3605 (.A(_04773_),
    .Y(net3605));
 BUFx3_ASAP7_75t_R place3606 (.A(_04770_),
    .Y(net3606));
 BUFx3_ASAP7_75t_R place3609 (.A(net3608),
    .Y(net3609));
 BUFx3_ASAP7_75t_R place3607 (.A(_03545_),
    .Y(net3607));
 BUFx3_ASAP7_75t_R place3608 (.A(_03534_),
    .Y(net3608));
 BUFx3_ASAP7_75t_R place3611 (.A(net3610),
    .Y(net3611));
 BUFx3_ASAP7_75t_R place3610 (.A(_03519_),
    .Y(net3610));
 BUFx6f_ASAP7_75t_R place3612 (.A(_03511_),
    .Y(net3612));
 BUFx3_ASAP7_75t_R place3614 (.A(_01845_),
    .Y(net3614));
 BUFx3_ASAP7_75t_R place3615 (.A(_01840_),
    .Y(net3615));
 BUFx3_ASAP7_75t_R place3616 (.A(_01819_),
    .Y(net3616));
 BUFx3_ASAP7_75t_R place3617 (.A(_01812_),
    .Y(net3617));
 BUFx3_ASAP7_75t_R place3619 (.A(_01799_),
    .Y(net3619));
 BUFx3_ASAP7_75t_R place3620 (.A(_05899_),
    .Y(net3620));
 BUFx3_ASAP7_75t_R place3621 (.A(_05894_),
    .Y(net3621));
 BUFx3_ASAP7_75t_R place3622 (.A(_05878_),
    .Y(net3622));
 BUFx3_ASAP7_75t_R place3624 (.A(net5611),
    .Y(net3624));
 BUFx3_ASAP7_75t_R place3625 (.A(_04820_),
    .Y(net3625));
 BUFx3_ASAP7_75t_R place3626 (.A(_04775_),
    .Y(net3626));
 BUFx3_ASAP7_75t_R place3627 (.A(_04772_),
    .Y(net3627));
 BUFx3_ASAP7_75t_R place3628 (.A(_04769_),
    .Y(net3628));
 BUFx3_ASAP7_75t_R place3629 (.A(_04764_),
    .Y(net3629));
 BUFx3_ASAP7_75t_R place3630 (.A(_04761_),
    .Y(net3630));
 BUFx3_ASAP7_75t_R place3631 (.A(_04750_),
    .Y(net3631));
 BUFx3_ASAP7_75t_R place3632 (.A(_03559_),
    .Y(net3632));
 BUFx3_ASAP7_75t_R place3634 (.A(_03549_),
    .Y(net3634));
 BUFx3_ASAP7_75t_R place3639 (.A(_01818_),
    .Y(net3639));
 BUFx3_ASAP7_75t_R place3637 (.A(_01823_),
    .Y(net3637));
 BUFx3_ASAP7_75t_R place3638 (.A(_01818_),
    .Y(net3638));
 BUFx3_ASAP7_75t_R place3640 (.A(_01811_),
    .Y(net3640));
 BUFx3_ASAP7_75t_R place3642 (.A(_01803_),
    .Y(net3642));
 BUFx3_ASAP7_75t_R place3643 (.A(_05870_),
    .Y(net3643));
 BUFx3_ASAP7_75t_R place3644 (.A(net5933),
    .Y(net3644));
 BUFx3_ASAP7_75t_R place3645 (.A(_04755_),
    .Y(net3645));
 BUFx3_ASAP7_75t_R place3647 (.A(_04736_),
    .Y(net3647));
 BUFx6f_ASAP7_75t_R rebuffer6002 (.A(_03411_),
    .Y(net6002));
 BUFx3_ASAP7_75t_R place3649 (.A(_03540_),
    .Y(net3649));
 BUFx3_ASAP7_75t_R place3656 (.A(_04733_),
    .Y(net3656));
 BUFx3_ASAP7_75t_R place3650 (.A(_03512_),
    .Y(net3650));
 BUFx3_ASAP7_75t_R place3651 (.A(_01801_),
    .Y(net3651));
 BUFx3_ASAP7_75t_R place3652 (.A(_01787_),
    .Y(net3652));
 BUFx3_ASAP7_75t_R place3655 (.A(_04748_),
    .Y(net3655));
 BUFx3_ASAP7_75t_R place3653 (.A(_04757_),
    .Y(net3653));
 BUFx3_ASAP7_75t_R place3654 (.A(_04748_),
    .Y(net3654));
 BUFx3_ASAP7_75t_R place3657 (.A(_04728_),
    .Y(net3657));
 BUFx3_ASAP7_75t_R place3658 (.A(_03538_),
    .Y(net3658));
 BUFx3_ASAP7_75t_R place3670 (.A(_04720_),
    .Y(net3670));
 BUFx3_ASAP7_75t_R place3660 (.A(_03514_),
    .Y(net3660));
 BUFx3_ASAP7_75t_R place3661 (.A(_03488_),
    .Y(net3661));
 BUFx3_ASAP7_75t_R place3662 (.A(_01814_),
    .Y(net3662));
 BUFx3_ASAP7_75t_R place3668 (.A(_04747_),
    .Y(net3668));
 BUFx3_ASAP7_75t_R place3663 (.A(_01786_),
    .Y(net3663));
 BUFx3_ASAP7_75t_R place3664 (.A(_05859_),
    .Y(net3664));
 BUFx3_ASAP7_75t_R place3665 (.A(_05847_),
    .Y(net3665));
 BUFx3_ASAP7_75t_R place3666 (.A(_04756_),
    .Y(net3666));
 BUFx3_ASAP7_75t_R place3667 (.A(_04754_),
    .Y(net3667));
 BUFx3_ASAP7_75t_R place3669 (.A(_04720_),
    .Y(net3669));
 BUFx3_ASAP7_75t_R place3671 (.A(_04709_),
    .Y(net3671));
 BUFx3_ASAP7_75t_R place3672 (.A(_03521_),
    .Y(net3672));
 BUFx3_ASAP7_75t_R place3673 (.A(_01800_),
    .Y(net3673));
 BUFx3_ASAP7_75t_R place3674 (.A(_01771_),
    .Y(net3674));
 BUFx3_ASAP7_75t_R place3675 (.A(_01765_),
    .Y(net3675));
 BUFx3_ASAP7_75t_R place3676 (.A(_01751_),
    .Y(net3676));
 BUFx3_ASAP7_75t_R place3681 (.A(_05825_),
    .Y(net3681));
 BUFx3_ASAP7_75t_R place3678 (.A(_05850_),
    .Y(net3678));
 BUFx3_ASAP7_75t_R place3679 (.A(_05842_),
    .Y(net3679));
 BUFx3_ASAP7_75t_R place3680 (.A(net5599),
    .Y(net3680));
 BUFx3_ASAP7_75t_R place3682 (.A(_05809_),
    .Y(net3682));
 BUFx3_ASAP7_75t_R place3683 (.A(_04746_),
    .Y(net3683));
 BUFx3_ASAP7_75t_R place3684 (.A(_04742_),
    .Y(net3684));
 BUFx3_ASAP7_75t_R place3703 (.A(_01795_),
    .Y(net3703));
 BUFx3_ASAP7_75t_R place3685 (.A(_04737_),
    .Y(net3685));
 BUFx3_ASAP7_75t_R place3686 (.A(_04732_),
    .Y(net3686));
 BUFx3_ASAP7_75t_R place3687 (.A(_04723_),
    .Y(net3687));
 BUFx3_ASAP7_75t_R place3702 (.A(_03486_),
    .Y(net3702));
 BUFx3_ASAP7_75t_R place3688 (.A(_04719_),
    .Y(net3688));
 BUFx3_ASAP7_75t_R place3694 (.A(_05817_),
    .Y(net3694));
 BUFx3_ASAP7_75t_R place3689 (.A(_04708_),
    .Y(net3689));
 BUFx3_ASAP7_75t_R place3690 (.A(_03509_),
    .Y(net3690));
 BUFx3_ASAP7_75t_R place3691 (.A(_01758_),
    .Y(net3691));
 BUFx3_ASAP7_75t_R place3692 (.A(_01750_),
    .Y(net3692));
 BUFx3_ASAP7_75t_R place3693 (.A(_05829_),
    .Y(net3693));
 BUFx3_ASAP7_75t_R place3695 (.A(_05808_),
    .Y(net3695));
 BUFx3_ASAP7_75t_R place3696 (.A(_04730_),
    .Y(net3696));
 BUFx3_ASAP7_75t_R place3697 (.A(_04729_),
    .Y(net3697));
 BUFx3_ASAP7_75t_R place3698 (.A(_04711_),
    .Y(net3698));
 BUFx3_ASAP7_75t_R place3699 (.A(_04707_),
    .Y(net3699));
 BUFx3_ASAP7_75t_R place3700 (.A(_04697_),
    .Y(net3700));
 BUFx3_ASAP7_75t_R place3701 (.A(_03490_),
    .Y(net3701));
 BUFx3_ASAP7_75t_R place3704 (.A(_01775_),
    .Y(net3704));
 BUFx3_ASAP7_75t_R place3706 (.A(_05851_),
    .Y(net3706));
 BUFx3_ASAP7_75t_R place3708 (.A(_05826_),
    .Y(net3708));
 BUFx3_ASAP7_75t_R place3709 (.A(_04696_),
    .Y(net3709));
 BUFx3_ASAP7_75t_R place3710 (.A(_03503_),
    .Y(net3710));
 BUFx3_ASAP7_75t_R place3712 (.A(_03485_),
    .Y(net3712));
 BUFx3_ASAP7_75t_R place3716 (.A(_05834_),
    .Y(net3716));
 BUFx3_ASAP7_75t_R place3717 (.A(_04738_),
    .Y(net3717));
 BUFx3_ASAP7_75t_R place3718 (.A(_04685_),
    .Y(net3718));
 BUFx3_ASAP7_75t_R place3723 (.A(_01762_),
    .Y(net3723));
 BUFx3_ASAP7_75t_R place3719 (.A(_03492_),
    .Y(net3719));
 BUFx3_ASAP7_75t_R place3720 (.A(_03489_),
    .Y(net3720));
 BUFx3_ASAP7_75t_R place3721 (.A(net5979),
    .Y(net3721));
 BUFx3_ASAP7_75t_R place3722 (.A(_01773_),
    .Y(net3722));
 BUFx3_ASAP7_75t_R place3724 (.A(_01747_),
    .Y(net3724));
 BUFx3_ASAP7_75t_R place3726 (.A(_01743_),
    .Y(net3726));
 BUFx3_ASAP7_75t_R place3729 (.A(net3728),
    .Y(net3729));
 BUFx3_ASAP7_75t_R place3728 (.A(_01738_),
    .Y(net3728));
 BUFx3_ASAP7_75t_R place3731 (.A(_01717_),
    .Y(net3731));
 BUFx3_ASAP7_75t_R place3730 (.A(_01717_),
    .Y(net3730));
 BUFx3_ASAP7_75t_R place3732 (.A(_05822_),
    .Y(net3732));
 BUFx3_ASAP7_75t_R place3733 (.A(_05804_),
    .Y(net3733));
 BUFx3_ASAP7_75t_R place3735 (.A(_05791_),
    .Y(net3735));
 BUFx3_ASAP7_75t_R place3736 (.A(_04731_),
    .Y(net3736));
 BUFx3_ASAP7_75t_R place3737 (.A(_04692_),
    .Y(net3737));
 BUFx3_ASAP7_75t_R place3738 (.A(_04684_),
    .Y(net3738));
 BUFx6f_ASAP7_75t_R place3739 (.A(_03447_),
    .Y(net3739));
 BUFx3_ASAP7_75t_R place3740 (.A(net5706),
    .Y(net3740));
 BUFx3_ASAP7_75t_R place3741 (.A(_01772_),
    .Y(net3741));
 BUFx3_ASAP7_75t_R place3742 (.A(_01766_),
    .Y(net3742));
 BUFx3_ASAP7_75t_R place3743 (.A(_01737_),
    .Y(net3743));
 BUFx3_ASAP7_75t_R place3744 (.A(_01734_),
    .Y(net3744));
 BUFx3_ASAP7_75t_R place3745 (.A(_01732_),
    .Y(net3745));
 BUFx3_ASAP7_75t_R place3746 (.A(net5763),
    .Y(net3746));
 BUFx3_ASAP7_75t_R place3747 (.A(_05797_),
    .Y(net3747));
 BUFx3_ASAP7_75t_R place3753 (.A(_03443_),
    .Y(net3753));
 BUFx3_ASAP7_75t_R place3748 (.A(_05777_),
    .Y(net3748));
 BUFx3_ASAP7_75t_R place3749 (.A(_05769_),
    .Y(net3749));
 BUFx3_ASAP7_75t_R place3750 (.A(_04714_),
    .Y(net3750));
 BUFx3_ASAP7_75t_R place3751 (.A(_04703_),
    .Y(net3751));
 BUFx3_ASAP7_75t_R place3752 (.A(_03483_),
    .Y(net3752));
 BUFx3_ASAP7_75t_R place3766 (.A(_04673_),
    .Y(net3766));
 BUFx3_ASAP7_75t_R place3764 (.A(_05765_),
    .Y(net3764));
 BUFx3_ASAP7_75t_R place3756 (.A(_04702_),
    .Y(net3756));
 BUFx3_ASAP7_75t_R place3757 (.A(_04698_),
    .Y(net3757));
 BUFx3_ASAP7_75t_R place3758 (.A(_04694_),
    .Y(net3758));
 BUFx3_ASAP7_75t_R place3759 (.A(_03453_),
    .Y(net3759));
 BUFx3_ASAP7_75t_R place3760 (.A(_01699_),
    .Y(net3760));
 BUFx3_ASAP7_75t_R place3761 (.A(_01684_),
    .Y(net3761));
 BUFx3_ASAP7_75t_R place3762 (.A(_05779_),
    .Y(net3762));
 BUFx3_ASAP7_75t_R place3763 (.A(_05767_),
    .Y(net3763));
 BUFx3_ASAP7_75t_R place3765 (.A(_04673_),
    .Y(net3765));
 BUFx3_ASAP7_75t_R place3767 (.A(net6010),
    .Y(net3767));
 BUFx3_ASAP7_75t_R place3768 (.A(_03441_),
    .Y(net3768));
 BUFx3_ASAP7_75t_R place3769 (.A(_03433_),
    .Y(net3769));
 BUFx3_ASAP7_75t_R place3774 (.A(net5771),
    .Y(net3774));
 BUFx3_ASAP7_75t_R place3771 (.A(_03424_),
    .Y(net3771));
 BUFx3_ASAP7_75t_R place3772 (.A(_01720_),
    .Y(net3772));
 BUFx3_ASAP7_75t_R place3773 (.A(_01714_),
    .Y(net3773));
 BUFx3_ASAP7_75t_R place3775 (.A(_01683_),
    .Y(net3775));
 BUFx3_ASAP7_75t_R place3782 (.A(net5617),
    .Y(net3782));
 BUFx3_ASAP7_75t_R place3778 (.A(_05784_),
    .Y(net3778));
 BUFx3_ASAP7_75t_R place3777 (.A(_05784_),
    .Y(net3777));
 BUFx3_ASAP7_75t_R place3779 (.A(_05778_),
    .Y(net3779));
 BUFx3_ASAP7_75t_R place3780 (.A(_05774_),
    .Y(net3780));
 BUFx6f_ASAP7_75t_R place3781 (.A(_05764_),
    .Y(net3781));
 BUFx3_ASAP7_75t_R place3783 (.A(_05731_),
    .Y(net3783));
 BUFx3_ASAP7_75t_R place3784 (.A(_04672_),
    .Y(net3784));
 BUFx3_ASAP7_75t_R place3785 (.A(_04663_),
    .Y(net3785));
 BUFx3_ASAP7_75t_R place3786 (.A(_04651_),
    .Y(net3786));
 BUFx3_ASAP7_75t_R place3787 (.A(_03445_),
    .Y(net3787));
 BUFx3_ASAP7_75t_R place3789 (.A(_03436_),
    .Y(net3789));
 BUFx3_ASAP7_75t_R place3791 (.A(net6002),
    .Y(net3791));
 BUFx3_ASAP7_75t_R place3792 (.A(_01703_),
    .Y(net3792));
 BUFx3_ASAP7_75t_R place3798 (.A(_05727_),
    .Y(net3798));
 BUFx3_ASAP7_75t_R place3794 (.A(_01682_),
    .Y(net3794));
 BUFx3_ASAP7_75t_R place3795 (.A(_01675_),
    .Y(net3795));
 BUFx3_ASAP7_75t_R place3796 (.A(net5961),
    .Y(net3796));
 BUFx3_ASAP7_75t_R place3797 (.A(_05757_),
    .Y(net3797));
 BUFx3_ASAP7_75t_R place3799 (.A(_04689_),
    .Y(net3799));
 BUFx3_ASAP7_75t_R place3800 (.A(_04678_),
    .Y(net3800));
 BUFx3_ASAP7_75t_R place3801 (.A(_04671_),
    .Y(net3801));
 BUFx3_ASAP7_75t_R place3802 (.A(_04650_),
    .Y(net3802));
 BUFx3_ASAP7_75t_R place3803 (.A(net5987),
    .Y(net3803));
 BUFx3_ASAP7_75t_R place3804 (.A(_03420_),
    .Y(net3804));
 BUFx6f_ASAP7_75t_R place3805 (.A(_01681_),
    .Y(net3805));
 BUFx3_ASAP7_75t_R place3806 (.A(_05762_),
    .Y(net3806));
 BUFx3_ASAP7_75t_R place3807 (.A(_05756_),
    .Y(net3807));
 BUFx3_ASAP7_75t_R place3809 (.A(_05726_),
    .Y(net3809));
 BUFx3_ASAP7_75t_R place3811 (.A(_04666_),
    .Y(net3811));
 BUFx3_ASAP7_75t_R place3813 (.A(_04655_),
    .Y(net3813));
 BUFx3_ASAP7_75t_R place3814 (.A(_04630_),
    .Y(net3814));
 BUFx3_ASAP7_75t_R place3815 (.A(_03417_),
    .Y(net3815));
 BUFx3_ASAP7_75t_R place3816 (.A(_03413_),
    .Y(net3816));
 BUFx3_ASAP7_75t_R place3817 (.A(_03409_),
    .Y(net3817));
 BUFx3_ASAP7_75t_R place3818 (.A(_01724_),
    .Y(net3818));
 BUFx3_ASAP7_75t_R place3819 (.A(_05761_),
    .Y(net3819));
 BUFx3_ASAP7_75t_R place3820 (.A(_05725_),
    .Y(net3820));
 BUFx3_ASAP7_75t_R place3824 (.A(_04634_),
    .Y(net3824));
 BUFx3_ASAP7_75t_R place3823 (.A(_04634_),
    .Y(net3823));
 BUFx3_ASAP7_75t_R place3825 (.A(_03412_),
    .Y(net3825));
 BUFx3_ASAP7_75t_R place3827 (.A(net6000),
    .Y(net3827));
 BUFx3_ASAP7_75t_R place3828 (.A(_03400_),
    .Y(net3828));
 BUFx3_ASAP7_75t_R place3829 (.A(_01696_),
    .Y(net3829));
 BUFx3_ASAP7_75t_R place3878 (.A(_03359_),
    .Y(net3878));
 BUFx3_ASAP7_75t_R place3830 (.A(_01690_),
    .Y(net3830));
 BUFx3_ASAP7_75t_R place3831 (.A(_01677_),
    .Y(net3831));
 BUFx3_ASAP7_75t_R place3832 (.A(_01676_),
    .Y(net3832));
 BUFx3_ASAP7_75t_R place3833 (.A(_01668_),
    .Y(net3833));
 BUFx3_ASAP7_75t_R place3841 (.A(_05701_),
    .Y(net3841));
 BUFx3_ASAP7_75t_R place3834 (.A(_05751_),
    .Y(net3834));
 BUFx3_ASAP7_75t_R place3835 (.A(_05747_),
    .Y(net3835));
 BUFx3_ASAP7_75t_R place3836 (.A(_05743_),
    .Y(net3836));
 BUFx3_ASAP7_75t_R place3837 (.A(_05738_),
    .Y(net3837));
 BUFx3_ASAP7_75t_R place3838 (.A(_05728_),
    .Y(net3838));
 BUFx3_ASAP7_75t_R place3839 (.A(_05713_),
    .Y(net3839));
 BUFx3_ASAP7_75t_R place3840 (.A(_05701_),
    .Y(net3840));
 BUFx3_ASAP7_75t_R place3848 (.A(net5697),
    .Y(net3848));
 BUFx3_ASAP7_75t_R place3842 (.A(_04654_),
    .Y(net3842));
 BUFx3_ASAP7_75t_R place3843 (.A(_04616_),
    .Y(net3843));
 BUFx3_ASAP7_75t_R place3844 (.A(_03406_),
    .Y(net3844));
 BUFx3_ASAP7_75t_R place3845 (.A(_03398_),
    .Y(net3845));
 BUFx3_ASAP7_75t_R place3846 (.A(_03389_),
    .Y(net3846));
 BUFx3_ASAP7_75t_R place3847 (.A(_03378_),
    .Y(net3847));
 BUFx3_ASAP7_75t_R place3858 (.A(_03401_),
    .Y(net3858));
 BUFx3_ASAP7_75t_R place3849 (.A(net5437),
    .Y(net3849));
 BUFx3_ASAP7_75t_R place3850 (.A(_05721_),
    .Y(net3850));
 BUFx3_ASAP7_75t_R place3851 (.A(_05700_),
    .Y(net3851));
 BUFx3_ASAP7_75t_R place3852 (.A(_04660_),
    .Y(net3852));
 BUFx3_ASAP7_75t_R place3853 (.A(_04647_),
    .Y(net3853));
 BUFx3_ASAP7_75t_R place3854 (.A(_04633_),
    .Y(net3854));
 BUFx3_ASAP7_75t_R place3855 (.A(_04629_),
    .Y(net3855));
 BUFx3_ASAP7_75t_R place3856 (.A(_04623_),
    .Y(net3856));
 BUFx3_ASAP7_75t_R place3857 (.A(_03405_),
    .Y(net3857));
 BUFx3_ASAP7_75t_R place3859 (.A(_03375_),
    .Y(net3859));
 BUFx3_ASAP7_75t_R place3860 (.A(_01673_),
    .Y(net3860));
 BUFx3_ASAP7_75t_R place3861 (.A(net5768),
    .Y(net3861));
 BUFx3_ASAP7_75t_R place3862 (.A(_01665_),
    .Y(net3862));
 BUFx3_ASAP7_75t_R place3863 (.A(_05735_),
    .Y(net3863));
 BUFx3_ASAP7_75t_R place3869 (.A(net5666),
    .Y(net3869));
 BUFx3_ASAP7_75t_R place3864 (.A(_05720_),
    .Y(net3864));
 BUFx3_ASAP7_75t_R place3865 (.A(_04637_),
    .Y(net3865));
 BUFx3_ASAP7_75t_R place3866 (.A(_04636_),
    .Y(net3866));
 BUFx3_ASAP7_75t_R place3867 (.A(_04604_),
    .Y(net3867));
 BUFx3_ASAP7_75t_R place3868 (.A(_04599_),
    .Y(net3868));
 BUFx3_ASAP7_75t_R place3870 (.A(_03374_),
    .Y(net3870));
 BUFx3_ASAP7_75t_R place3871 (.A(_01654_),
    .Y(net3871));
 BUFx3_ASAP7_75t_R place3872 (.A(_05734_),
    .Y(net3872));
 BUFx3_ASAP7_75t_R place3873 (.A(_04613_),
    .Y(net3873));
 BUFx3_ASAP7_75t_R place3874 (.A(_04611_),
    .Y(net3874));
 BUFx3_ASAP7_75t_R place3875 (.A(_04600_),
    .Y(net3875));
 BUFx3_ASAP7_75t_R place3876 (.A(_03373_),
    .Y(net3876));
 BUFx3_ASAP7_75t_R place3877 (.A(_03359_),
    .Y(net3877));
 BUFx3_ASAP7_75t_R place3881 (.A(net3880),
    .Y(net3881));
 BUFx3_ASAP7_75t_R place3879 (.A(_05723_),
    .Y(net3879));
 BUFx3_ASAP7_75t_R place3880 (.A(_05710_),
    .Y(net3880));
 BUFx3_ASAP7_75t_R place3913 (.A(net3912),
    .Y(net3913));
 BUFx3_ASAP7_75t_R place3882 (.A(_05708_),
    .Y(net3882));
 BUFx3_ASAP7_75t_R place3883 (.A(_05705_),
    .Y(net3883));
 BUFx6f_ASAP7_75t_R place3884 (.A(_05670_),
    .Y(net3884));
 BUFx3_ASAP7_75t_R place3889 (.A(_03372_),
    .Y(net3889));
 BUFx3_ASAP7_75t_R place3885 (.A(_04587_),
    .Y(net3885));
 BUFx3_ASAP7_75t_R place3886 (.A(_04565_),
    .Y(net3886));
 BUFx3_ASAP7_75t_R place3887 (.A(_03404_),
    .Y(net3887));
 BUFx3_ASAP7_75t_R place3888 (.A(_03380_),
    .Y(net3888));
 BUFx3_ASAP7_75t_R place3890 (.A(net5977),
    .Y(net3890));
 BUFx3_ASAP7_75t_R place3891 (.A(_01657_),
    .Y(net3891));
 BUFx3_ASAP7_75t_R place3892 (.A(_01635_),
    .Y(net3892));
 BUFx3_ASAP7_75t_R place3893 (.A(_01630_),
    .Y(net3893));
 BUFx3_ASAP7_75t_R place3894 (.A(_01609_),
    .Y(net3894));
 BUFx3_ASAP7_75t_R place3895 (.A(_05698_),
    .Y(net3895));
 BUFx3_ASAP7_75t_R place3896 (.A(_05693_),
    .Y(net3896));
 BUFx3_ASAP7_75t_R place3897 (.A(_04607_),
    .Y(net3897));
 BUFx3_ASAP7_75t_R place3901 (.A(_04586_),
    .Y(net3901));
 BUFx3_ASAP7_75t_R place3898 (.A(_04603_),
    .Y(net3898));
 BUFx3_ASAP7_75t_R place3899 (.A(_04596_),
    .Y(net3899));
 BUFx3_ASAP7_75t_R place3900 (.A(_04588_),
    .Y(net3900));
 BUFx3_ASAP7_75t_R place3902 (.A(_03395_),
    .Y(net3902));
 BUFx3_ASAP7_75t_R place3903 (.A(_03370_),
    .Y(net3903));
 BUFx3_ASAP7_75t_R place3904 (.A(_03364_),
    .Y(net3904));
 BUFx3_ASAP7_75t_R place3905 (.A(_01655_),
    .Y(net3905));
 BUFx3_ASAP7_75t_R place3906 (.A(_01643_),
    .Y(net3906));
 BUFx3_ASAP7_75t_R place3907 (.A(_05680_),
    .Y(net3907));
 BUFx3_ASAP7_75t_R place3908 (.A(net5938),
    .Y(net3908));
 BUFx3_ASAP7_75t_R place3909 (.A(_04617_),
    .Y(net3909));
 BUFx3_ASAP7_75t_R place3910 (.A(_04563_),
    .Y(net3910));
 BUFx3_ASAP7_75t_R place3912 (.A(_03368_),
    .Y(net3912));
 BUFx3_ASAP7_75t_R place3911 (.A(_03369_),
    .Y(net3911));
 BUFx3_ASAP7_75t_R place3914 (.A(_03351_),
    .Y(net3914));
 BUFx3_ASAP7_75t_R place3915 (.A(_01628_),
    .Y(net3915));
 BUFx3_ASAP7_75t_R place3916 (.A(_05690_),
    .Y(net3916));
 BUFx3_ASAP7_75t_R place3920 (.A(_04560_),
    .Y(net3920));
 BUFx3_ASAP7_75t_R place3917 (.A(_05679_),
    .Y(net3917));
 BUFx3_ASAP7_75t_R place3918 (.A(_04570_),
    .Y(net3918));
 BUFx6f_ASAP7_75t_R place3919 (.A(_04569_),
    .Y(net3919));
 BUFx3_ASAP7_75t_R place3921 (.A(net5680),
    .Y(net3921));
 BUFx3_ASAP7_75t_R place3923 (.A(_01620_),
    .Y(net3923));
 BUFx3_ASAP7_75t_R place3924 (.A(_01618_),
    .Y(net3924));
 BUFx3_ASAP7_75t_R place3925 (.A(_01616_),
    .Y(net3925));
 BUFx3_ASAP7_75t_R place3926 (.A(_01605_),
    .Y(net3926));
 BUFx3_ASAP7_75t_R place3928 (.A(_05672_),
    .Y(net3928));
 BUFx3_ASAP7_75t_R place3929 (.A(_05665_),
    .Y(net3929));
 BUFx3_ASAP7_75t_R place3930 (.A(_04559_),
    .Y(net3930));
 BUFx3_ASAP7_75t_R place3932 (.A(_04557_),
    .Y(net3932));
 BUFx3_ASAP7_75t_R place3933 (.A(_04539_),
    .Y(net3933));
 BUFx3_ASAP7_75t_R place3935 (.A(_01603_),
    .Y(net3935));
 BUFx3_ASAP7_75t_R place3939 (.A(net3938),
    .Y(net3939));
 BUFx3_ASAP7_75t_R place3936 (.A(net5430),
    .Y(net3936));
 BUFx3_ASAP7_75t_R place3937 (.A(_05671_),
    .Y(net3937));
 BUFx6f_ASAP7_75t_R place3938 (.A(_05636_),
    .Y(net3938));
 BUFx3_ASAP7_75t_R place3941 (.A(_04558_),
    .Y(net3941));
 BUFx3_ASAP7_75t_R place3942 (.A(_04543_),
    .Y(net3942));
 BUFx3_ASAP7_75t_R place3943 (.A(_04538_),
    .Y(net3943));
 BUFx6f_ASAP7_75t_R place3944 (.A(_03367_),
    .Y(net3944));
 BUFx3_ASAP7_75t_R place3945 (.A(_03348_),
    .Y(net3945));
 BUFx3_ASAP7_75t_R place3946 (.A(_05664_),
    .Y(net3946));
 BUFx3_ASAP7_75t_R place3947 (.A(_05639_),
    .Y(net3947));
 BUFx3_ASAP7_75t_R place3948 (.A(_04578_),
    .Y(net3948));
 BUFx3_ASAP7_75t_R place3949 (.A(_04550_),
    .Y(net3949));
 BUFx3_ASAP7_75t_R place3950 (.A(_04541_),
    .Y(net3950));
 BUFx3_ASAP7_75t_R place3951 (.A(_03347_),
    .Y(net3951));
 BUFx3_ASAP7_75t_R place3952 (.A(_01592_),
    .Y(net3952));
 BUFx3_ASAP7_75t_R place3954 (.A(net5959),
    .Y(net3954));
 BUFx3_ASAP7_75t_R place3955 (.A(_05642_),
    .Y(net3955));
 BUFx3_ASAP7_75t_R place3956 (.A(_05638_),
    .Y(net3956));
 BUFx3_ASAP7_75t_R place3979 (.A(_04542_),
    .Y(net3979));
 BUFx3_ASAP7_75t_R place3957 (.A(_05597_),
    .Y(net3957));
 BUFx3_ASAP7_75t_R place3958 (.A(_04576_),
    .Y(net3958));
 BUFx3_ASAP7_75t_R place3959 (.A(_04548_),
    .Y(net3959));
 BUFx3_ASAP7_75t_R place3960 (.A(_04529_),
    .Y(net3960));
 BUFx3_ASAP7_75t_R place3965 (.A(_01549_),
    .Y(net3965));
 BUFx3_ASAP7_75t_R place3961 (.A(_03353_),
    .Y(net3961));
 BUFx3_ASAP7_75t_R place3962 (.A(_03337_),
    .Y(net3962));
 BUFx3_ASAP7_75t_R place3963 (.A(_01589_),
    .Y(net3963));
 BUFx3_ASAP7_75t_R place3964 (.A(_01549_),
    .Y(net3964));
 BUFx3_ASAP7_75t_R place3974 (.A(_01520_),
    .Y(net3974));
 BUFx3_ASAP7_75t_R place3966 (.A(_05634_),
    .Y(net3966));
 BUFx3_ASAP7_75t_R place3967 (.A(_05607_),
    .Y(net3967));
 BUFx3_ASAP7_75t_R place3968 (.A(_05596_),
    .Y(net3968));
 BUFx3_ASAP7_75t_R place3969 (.A(_04536_),
    .Y(net3969));
 BUFx3_ASAP7_75t_R place3973 (.A(_01520_),
    .Y(net3973));
 BUFx3_ASAP7_75t_R place3970 (.A(_03339_),
    .Y(net3970));
 BUFx3_ASAP7_75t_R place3971 (.A(_01548_),
    .Y(net3971));
 BUFx3_ASAP7_75t_R place3972 (.A(_01527_),
    .Y(net3972));
 BUFx3_ASAP7_75t_R place3975 (.A(_01515_),
    .Y(net3975));
 BUFx3_ASAP7_75t_R place3976 (.A(_05606_),
    .Y(net3976));
 BUFx3_ASAP7_75t_R place3977 (.A(_04547_),
    .Y(net3977));
 BUFx3_ASAP7_75t_R place3978 (.A(_04544_),
    .Y(net3978));
 BUFx3_ASAP7_75t_R place3980 (.A(_04533_),
    .Y(net3980));
 BUFx3_ASAP7_75t_R place3981 (.A(_04505_),
    .Y(net3981));
 BUFx3_ASAP7_75t_R place3982 (.A(_03334_),
    .Y(net3982));
 BUFx3_ASAP7_75t_R place3985 (.A(_01519_),
    .Y(net3985));
 BUFx3_ASAP7_75t_R place3986 (.A(_04532_),
    .Y(net3986));
 BUFx3_ASAP7_75t_R place3987 (.A(_04504_),
    .Y(net3987));
 BUFx3_ASAP7_75t_R place3989 (.A(net5716),
    .Y(net3989));
 BUFx3_ASAP7_75t_R place3990 (.A(_01533_),
    .Y(net3990));
 BUFx3_ASAP7_75t_R place3991 (.A(_01532_),
    .Y(net3991));
 BUFx3_ASAP7_75t_R place4028 (.A(_05810_),
    .Y(net4028));
 BUFx6f_ASAP7_75t_R place3992 (.A(_05631_),
    .Y(net3992));
 BUFx3_ASAP7_75t_R place4021 (.A(_02809_),
    .Y(net4021));
 BUFx3_ASAP7_75t_R place3993 (.A(_04556_),
    .Y(net3993));
 BUFx3_ASAP7_75t_R place3994 (.A(_04535_),
    .Y(net3994));
 BUFx6f_ASAP7_75t_R place3999 (.A(_02899_),
    .Y(net3999));
 BUFx3_ASAP7_75t_R place3995 (.A(_04486_),
    .Y(net3995));
 BUFx3_ASAP7_75t_R place3996 (.A(_03328_),
    .Y(net3996));
 BUFx3_ASAP7_75t_R place3997 (.A(_03307_),
    .Y(net3997));
 BUFx6f_ASAP7_75t_R place3998 (.A(_02899_),
    .Y(net3998));
 BUFx3_ASAP7_75t_R place4020 (.A(_02809_),
    .Y(net4020));
 BUFx3_ASAP7_75t_R place4000 (.A(net6030),
    .Y(net4000));
 BUFx12f_ASAP7_75t_R place4018 (.A(net4015),
    .Y(net4018));
 BUFx12f_ASAP7_75t_R place4016 (.A(net4015),
    .Y(net4016));
 BUFx3_ASAP7_75t_R place4008 (.A(net4007),
    .Y(net4008));
 BUFx3_ASAP7_75t_R place4004 (.A(_05663_),
    .Y(net4004));
 BUFx6f_ASAP7_75t_R place4017 (.A(net4015),
    .Y(net4017));
 BUFx3_ASAP7_75t_R place4001 (.A(_01512_),
    .Y(net4001));
 BUFx3_ASAP7_75t_R place4002 (.A(_01469_),
    .Y(net4002));
 BUFx6f_ASAP7_75t_R place4003 (.A(_05663_),
    .Y(net4003));
 BUFx3_ASAP7_75t_R place4005 (.A(_05592_),
    .Y(net4005));
 BUFx3_ASAP7_75t_R place4006 (.A(_04555_),
    .Y(net4006));
 BUFx3_ASAP7_75t_R place4007 (.A(_04528_),
    .Y(net4007));
 BUFx3_ASAP7_75t_R place4010 (.A(_04503_),
    .Y(net4010));
 BUFx3_ASAP7_75t_R place4009 (.A(_04525_),
    .Y(net4009));
 BUFx3_ASAP7_75t_R place4011 (.A(_04468_),
    .Y(net4011));
 BUFx3_ASAP7_75t_R place4012 (.A(_03327_),
    .Y(net4012));
 BUFx3_ASAP7_75t_R place4013 (.A(_03325_),
    .Y(net4013));
 BUFx3_ASAP7_75t_R place4014 (.A(_03297_),
    .Y(net4014));
 BUFx6f_ASAP7_75t_R place4015 (.A(_02897_),
    .Y(net4015));
 BUFx3_ASAP7_75t_R place4019 (.A(net6041),
    .Y(net4019));
 BUFx3_ASAP7_75t_R place4022 (.A(_02367_),
    .Y(net4022));
 BUFx3_ASAP7_75t_R place4023 (.A(_01782_),
    .Y(net4023));
 BUFx3_ASAP7_75t_R place4024 (.A(_01656_),
    .Y(net4024));
 BUFx3_ASAP7_75t_R place4025 (.A(_01559_),
    .Y(net4025));
 BUFx3_ASAP7_75t_R place4026 (.A(_01468_),
    .Y(net4026));
 BUFx3_ASAP7_75t_R place4027 (.A(_05810_),
    .Y(net4027));
 BUFx3_ASAP7_75t_R place4029 (.A(_05749_),
    .Y(net4029));
 BUFx3_ASAP7_75t_R place4030 (.A(_05662_),
    .Y(net4030));
 BUFx3_ASAP7_75t_R place4031 (.A(_05637_),
    .Y(net4031));
 BUFx3_ASAP7_75t_R place4032 (.A(_05617_),
    .Y(net4032));
 BUFx3_ASAP7_75t_R place4037 (.A(_04467_),
    .Y(net4037));
 BUFx3_ASAP7_75t_R place4033 (.A(_04638_),
    .Y(net4033));
 BUFx3_ASAP7_75t_R place4034 (.A(_04621_),
    .Y(net4034));
 BUFx3_ASAP7_75t_R place4035 (.A(_04527_),
    .Y(net4035));
 BUFx3_ASAP7_75t_R place4036 (.A(_04502_),
    .Y(net4036));
 BUFx3_ASAP7_75t_R place4038 (.A(_03516_),
    .Y(net4038));
 BUFx3_ASAP7_75t_R place4039 (.A(_03440_),
    .Y(net4039));
 BUFx3_ASAP7_75t_R place4040 (.A(_03302_),
    .Y(net4040));
 BUFx6f_ASAP7_75t_R place4043 (.A(net6038),
    .Y(net4043));
 BUFx3_ASAP7_75t_R place4042 (.A(_02975_),
    .Y(net4042));
 BUFx3_ASAP7_75t_R place4044 (.A(_02811_),
    .Y(net4044));
 BUFx3_ASAP7_75t_R place4045 (.A(_02807_),
    .Y(net4045));
 BUFx3_ASAP7_75t_R place4046 (.A(_02364_),
    .Y(net4046));
 BUFx3_ASAP7_75t_R place4047 (.A(_01834_),
    .Y(net4047));
 BUFx3_ASAP7_75t_R place4048 (.A(_01761_),
    .Y(net4048));
 BUFx3_ASAP7_75t_R place4049 (.A(_01695_),
    .Y(net4049));
 BUFx3_ASAP7_75t_R place4050 (.A(_01642_),
    .Y(net4050));
 BUFx6f_ASAP7_75t_R place4051 (.A(_01557_),
    .Y(net4051));
 BUFx3_ASAP7_75t_R place4064 (.A(net4063),
    .Y(net4064));
 BUFx3_ASAP7_75t_R place4053 (.A(_01524_),
    .Y(net4053));
 BUFx3_ASAP7_75t_R place4054 (.A(_01498_),
    .Y(net4054));
 BUFx3_ASAP7_75t_R place4055 (.A(_01486_),
    .Y(net4055));
 BUFx3_ASAP7_75t_R place4056 (.A(net5425),
    .Y(net4056));
 BUFx3_ASAP7_75t_R place4057 (.A(_05918_),
    .Y(net4057));
 BUFx3_ASAP7_75t_R place4061 (.A(net4060),
    .Y(net4061));
 BUFx3_ASAP7_75t_R place4058 (.A(_05871_),
    .Y(net4058));
 BUFx3_ASAP7_75t_R place4059 (.A(_05800_),
    .Y(net4059));
 BUFx3_ASAP7_75t_R place4060 (.A(_05716_),
    .Y(net4060));
 BUFx3_ASAP7_75t_R place4062 (.A(_05683_),
    .Y(net4062));
 BUFx3_ASAP7_75t_R place4063 (.A(_05620_),
    .Y(net4063));
 BUFx3_ASAP7_75t_R place4066 (.A(_04823_),
    .Y(net4066));
 BUFx3_ASAP7_75t_R place4067 (.A(_04768_),
    .Y(net4067));
 BUFx3_ASAP7_75t_R place4068 (.A(_04727_),
    .Y(net4068));
 BUFx3_ASAP7_75t_R place4070 (.A(_04620_),
    .Y(net4070));
 BUFx3_ASAP7_75t_R place4071 (.A(_04562_),
    .Y(net4071));
 BUFx3_ASAP7_75t_R place4072 (.A(_04491_),
    .Y(net4072));
 BUFx3_ASAP7_75t_R place4073 (.A(_04422_),
    .Y(net4073));
 BUFx3_ASAP7_75t_R place4074 (.A(_03750_),
    .Y(net4074));
 BUFx3_ASAP7_75t_R place4084 (.A(_03264_),
    .Y(net4084));
 BUFx3_ASAP7_75t_R place4076 (.A(_03698_),
    .Y(net4076));
 BUFx3_ASAP7_75t_R place4077 (.A(_03631_),
    .Y(net4077));
 BUFx3_ASAP7_75t_R place4078 (.A(_03568_),
    .Y(net4078));
 BUFx3_ASAP7_75t_R place4079 (.A(_03496_),
    .Y(net4079));
 BUFx3_ASAP7_75t_R place4080 (.A(_03423_),
    .Y(net4080));
 BUFx3_ASAP7_75t_R place4081 (.A(_03407_),
    .Y(net4081));
 BUFx3_ASAP7_75t_R place4082 (.A(_03371_),
    .Y(net4082));
 BUFx3_ASAP7_75t_R place4083 (.A(_03324_),
    .Y(net4083));
 BUFx6f_ASAP7_75t_R place4085 (.A(net6027),
    .Y(net4085));
 BUFx6f_ASAP7_75t_R place4087 (.A(_02806_),
    .Y(net4087));
 BUFx3_ASAP7_75t_R place4088 (.A(_02378_),
    .Y(net4088));
 BUFx3_ASAP7_75t_R place4089 (.A(_02311_),
    .Y(net4089));
 BUFx3_ASAP7_75t_R place4090 (.A(_02249_),
    .Y(net4090));
 BUFx3_ASAP7_75t_R place4091 (.A(_02156_),
    .Y(net4091));
 BUFx3_ASAP7_75t_R place4092 (.A(_02137_),
    .Y(net4092));
 BUFx3_ASAP7_75t_R place4093 (.A(_01938_),
    .Y(net4093));
 BUFx6f_ASAP7_75t_R place4094 (.A(_01934_),
    .Y(net4094));
 BUFx3_ASAP7_75t_R place4095 (.A(_01857_),
    .Y(net4095));
 BUFx3_ASAP7_75t_R place4096 (.A(_01833_),
    .Y(net4096));
 BUFx3_ASAP7_75t_R place4097 (.A(_01817_),
    .Y(net4097));
 BUFx3_ASAP7_75t_R place4098 (.A(_01710_),
    .Y(net4098));
 BUFx3_ASAP7_75t_R place4099 (.A(_01686_),
    .Y(net4099));
 BUFx3_ASAP7_75t_R place4100 (.A(_01600_),
    .Y(net4100));
 BUFx3_ASAP7_75t_R place4101 (.A(_01334_),
    .Y(net4101));
 BUFx3_ASAP7_75t_R place4102 (.A(_01179_),
    .Y(net4102));
 BUFx3_ASAP7_75t_R place4103 (.A(_01163_),
    .Y(net4103));
 BUFx6f_ASAP7_75t_R place4104 (.A(net5730),
    .Y(net4104));
 BUFx3_ASAP7_75t_R place4105 (.A(_06504_),
    .Y(net4105));
 BUFx3_ASAP7_75t_R place4108 (.A(_05908_),
    .Y(net4108));
 BUFx3_ASAP7_75t_R place4110 (.A(net4109),
    .Y(net4110));
 BUFx3_ASAP7_75t_R place4109 (.A(_05865_),
    .Y(net4109));
 BUFx3_ASAP7_75t_R place4114 (.A(net4113),
    .Y(net4114));
 BUFx3_ASAP7_75t_R place4111 (.A(_05832_),
    .Y(net4111));
 BUFx3_ASAP7_75t_R place4112 (.A(_05682_),
    .Y(net4112));
 BUFx3_ASAP7_75t_R place4113 (.A(_05210_),
    .Y(net4113));
 BUFx3_ASAP7_75t_R place4122 (.A(_04895_),
    .Y(net4122));
 BUFx3_ASAP7_75t_R place4115 (.A(_05139_),
    .Y(net4115));
 BUFx3_ASAP7_75t_R place4116 (.A(_05121_),
    .Y(net4116));
 BUFx3_ASAP7_75t_R place4117 (.A(_05072_),
    .Y(net4117));
 BUFx3_ASAP7_75t_R place4118 (.A(_04987_),
    .Y(net4118));
 BUFx3_ASAP7_75t_R place4119 (.A(_04945_),
    .Y(net4119));
 BUFx3_ASAP7_75t_R place4120 (.A(_04906_),
    .Y(net4120));
 BUFx3_ASAP7_75t_R place4121 (.A(_04895_),
    .Y(net4121));
 BUFx3_ASAP7_75t_R place4123 (.A(_04836_),
    .Y(net4123));
 BUFx6f_ASAP7_75t_R place4124 (.A(_04790_),
    .Y(net4124));
 BUFx3_ASAP7_75t_R place4126 (.A(_04735_),
    .Y(net4126));
 BUFx3_ASAP7_75t_R place4127 (.A(_04726_),
    .Y(net4127));
 BUFx3_ASAP7_75t_R place4130 (.A(net4129),
    .Y(net4130));
 BUFx3_ASAP7_75t_R place4129 (.A(_04657_),
    .Y(net4129));
 BUFx3_ASAP7_75t_R place4131 (.A(_04497_),
    .Y(net4131));
 BUFx3_ASAP7_75t_R place4132 (.A(_04421_),
    .Y(net4132));
 BUFx3_ASAP7_75t_R place4134 (.A(_04092_),
    .Y(net4134));
 BUFx3_ASAP7_75t_R place4136 (.A(_03984_),
    .Y(net4136));
 BUFx6f_ASAP7_75t_R place4135 (.A(_04041_),
    .Y(net4135));
 BUFx3_ASAP7_75t_R place4143 (.A(net4142),
    .Y(net4143));
 BUFx3_ASAP7_75t_R place4137 (.A(_03906_),
    .Y(net4137));
 BUFx3_ASAP7_75t_R place4138 (.A(_03785_),
    .Y(net4138));
 BUFx3_ASAP7_75t_R place4139 (.A(_03749_),
    .Y(net4139));
 BUFx3_ASAP7_75t_R place4140 (.A(_03744_),
    .Y(net4140));
 BUFx3_ASAP7_75t_R place4141 (.A(_03678_),
    .Y(net4141));
 BUFx6f_ASAP7_75t_R place4142 (.A(_03630_),
    .Y(net4142));
 BUFx3_ASAP7_75t_R place4144 (.A(_03567_),
    .Y(net4144));
 BUFx3_ASAP7_75t_R place4145 (.A(_03462_),
    .Y(net4145));
 BUFx6f_ASAP7_75t_R place4146 (.A(_03388_),
    .Y(net4146));
 BUFx3_ASAP7_75t_R place4148 (.A(_03323_),
    .Y(net4148));
 BUFx3_ASAP7_75t_R place4149 (.A(_03314_),
    .Y(net4149));
 BUFx3_ASAP7_75t_R place4150 (.A(_03287_),
    .Y(net4150));
 BUFx3_ASAP7_75t_R place4151 (.A(net6042),
    .Y(net4151));
 BUFx3_ASAP7_75t_R place4152 (.A(_01100_),
    .Y(net4152));
 BUFx3_ASAP7_75t_R place4153 (.A(_02363_),
    .Y(net4153));
 BUFx3_ASAP7_75t_R place4154 (.A(_02310_),
    .Y(net4154));
 BUFx3_ASAP7_75t_R place4155 (.A(_02248_),
    .Y(net4155));
 BUFx3_ASAP7_75t_R place4156 (.A(_02168_),
    .Y(net4156));
 BUFx3_ASAP7_75t_R place4158 (.A(_02155_),
    .Y(net4158));
 BUFx3_ASAP7_75t_R place4159 (.A(_02107_),
    .Y(net4159));
 BUFx3_ASAP7_75t_R place4161 (.A(_02088_),
    .Y(net4161));
 BUFx3_ASAP7_75t_R place4164 (.A(_01985_),
    .Y(net4164));
 BUFx3_ASAP7_75t_R place4165 (.A(_01937_),
    .Y(net4165));
 BUFx3_ASAP7_75t_R place4166 (.A(_01911_),
    .Y(net4166));
 BUFx3_ASAP7_75t_R place4168 (.A(_01856_),
    .Y(net4168));
 BUFx3_ASAP7_75t_R place4171 (.A(net4170),
    .Y(net4171));
 BUFx3_ASAP7_75t_R place4170 (.A(_01806_),
    .Y(net4170));
 BUFx3_ASAP7_75t_R place4172 (.A(_01709_),
    .Y(net4172));
 BUFx3_ASAP7_75t_R place4173 (.A(_01640_),
    .Y(net4173));
 BUFx3_ASAP7_75t_R place4174 (.A(_01564_),
    .Y(net4174));
 BUFx3_ASAP7_75t_R place4175 (.A(_01488_),
    .Y(net4175));
 BUFx3_ASAP7_75t_R place4176 (.A(_01333_),
    .Y(net4176));
 BUFx3_ASAP7_75t_R place4177 (.A(_01178_),
    .Y(net4177));
 BUFx3_ASAP7_75t_R place4178 (.A(_01162_),
    .Y(net4178));
 BUFx3_ASAP7_75t_R place4179 (.A(_01119_),
    .Y(net4179));
 BUFx3_ASAP7_75t_R place4180 (.A(_06095_),
    .Y(net4180));
 BUFx3_ASAP7_75t_R place4189 (.A(net4188),
    .Y(net4189));
 BUFx3_ASAP7_75t_R place4182 (.A(_06006_),
    .Y(net4182));
 BUFx3_ASAP7_75t_R place4183 (.A(_05978_),
    .Y(net4183));
 BUFx3_ASAP7_75t_R place4184 (.A(_05889_),
    .Y(net4184));
 BUFx3_ASAP7_75t_R place4185 (.A(_05831_),
    .Y(net4185));
 BUFx3_ASAP7_75t_R place4186 (.A(_05759_),
    .Y(net4186));
 BUFx3_ASAP7_75t_R place4187 (.A(_05659_),
    .Y(net4187));
 BUFx3_ASAP7_75t_R place4188 (.A(_05602_),
    .Y(net4188));
 BUFx3_ASAP7_75t_R place4190 (.A(_05549_),
    .Y(net4190));
 BUFx3_ASAP7_75t_R place4191 (.A(_05351_),
    .Y(net4191));
 BUFx3_ASAP7_75t_R place4192 (.A(_05209_),
    .Y(net4192));
 BUFx3_ASAP7_75t_R place4193 (.A(_05138_),
    .Y(net4193));
 BUFx3_ASAP7_75t_R place4194 (.A(_05100_),
    .Y(net4194));
 BUFx3_ASAP7_75t_R place4196 (.A(_05060_),
    .Y(net4196));
 BUFx3_ASAP7_75t_R place4195 (.A(_05060_),
    .Y(net4195));
 BUFx3_ASAP7_75t_R place4210 (.A(_04066_),
    .Y(net4210));
 BUFx3_ASAP7_75t_R place4197 (.A(_05011_),
    .Y(net4197));
 BUFx3_ASAP7_75t_R place4198 (.A(_04986_),
    .Y(net4198));
 BUFx3_ASAP7_75t_R place4199 (.A(_04944_),
    .Y(net4199));
 BUFx3_ASAP7_75t_R place4200 (.A(_04905_),
    .Y(net4200));
 BUFx3_ASAP7_75t_R place4201 (.A(_04868_),
    .Y(net4201));
 BUFx3_ASAP7_75t_R place4207 (.A(_04368_),
    .Y(net4207));
 BUFx6f_ASAP7_75t_R place4203 (.A(_04835_),
    .Y(net4203));
 BUFx3_ASAP7_75t_R place4202 (.A(_04835_),
    .Y(net4202));
 BUFx3_ASAP7_75t_R place4204 (.A(_04495_),
    .Y(net4204));
 BUFx3_ASAP7_75t_R place4205 (.A(_04465_),
    .Y(net4205));
 BUFx3_ASAP7_75t_R place4206 (.A(_04459_),
    .Y(net4206));
 BUFx3_ASAP7_75t_R place4208 (.A(_04111_),
    .Y(net4208));
 BUFx3_ASAP7_75t_R place4209 (.A(_04066_),
    .Y(net4209));
 BUFx3_ASAP7_75t_R place4211 (.A(_03999_),
    .Y(net4211));
 BUFx3_ASAP7_75t_R place4212 (.A(_03973_),
    .Y(net4212));
 BUFx3_ASAP7_75t_R place4246 (.A(net4245),
    .Y(net4246));
 BUFx3_ASAP7_75t_R place4213 (.A(_03921_),
    .Y(net4213));
 BUFx3_ASAP7_75t_R place4214 (.A(_03905_),
    .Y(net4214));
 BUFx3_ASAP7_75t_R place4236 (.A(_01081_),
    .Y(net4236));
 BUFx3_ASAP7_75t_R place4215 (.A(_03784_),
    .Y(net4215));
 BUFx3_ASAP7_75t_R place4216 (.A(_03705_),
    .Y(net4216));
 BUFx3_ASAP7_75t_R place4217 (.A(_03612_),
    .Y(net4217));
 BUFx3_ASAP7_75t_R place4228 (.A(net4227),
    .Y(net4228));
 BUFx3_ASAP7_75t_R place4218 (.A(_03561_),
    .Y(net4218));
 BUFx3_ASAP7_75t_R place4219 (.A(_03247_),
    .Y(net4219));
 BUFx3_ASAP7_75t_R place4220 (.A(_03186_),
    .Y(net4220));
 BUFx3_ASAP7_75t_R place4221 (.A(_03170_),
    .Y(net4221));
 BUFx3_ASAP7_75t_R place4222 (.A(_02769_),
    .Y(net4222));
 BUFx3_ASAP7_75t_R place4223 (.A(_02639_),
    .Y(net4223));
 BUFx3_ASAP7_75t_R place4224 (.A(_01099_),
    .Y(net4224));
 BUFx3_ASAP7_75t_R place4225 (.A(_02366_),
    .Y(net4225));
 BUFx3_ASAP7_75t_R place4226 (.A(_02167_),
    .Y(net4226));
 BUFx3_ASAP7_75t_R place4227 (.A(_02036_),
    .Y(net4227));
 BUFx3_ASAP7_75t_R place4229 (.A(_01577_),
    .Y(net4229));
 BUFx3_ASAP7_75t_R place4230 (.A(_01544_),
    .Y(net4230));
 BUFx3_ASAP7_75t_R place4231 (.A(_01542_),
    .Y(net4231));
 BUFx3_ASAP7_75t_R place4232 (.A(_01541_),
    .Y(net4232));
 BUFx3_ASAP7_75t_R place4233 (.A(_01487_),
    .Y(net4233));
 BUFx3_ASAP7_75t_R place4234 (.A(_01452_),
    .Y(net4234));
 BUFx3_ASAP7_75t_R place4235 (.A(_01118_),
    .Y(net4235));
 BUFx3_ASAP7_75t_R place4237 (.A(_06373_),
    .Y(net4237));
 BUFx3_ASAP7_75t_R place4238 (.A(_06367_),
    .Y(net4238));
 BUFx3_ASAP7_75t_R place4239 (.A(_06312_),
    .Y(net4239));
 BUFx6f_ASAP7_75t_R place4240 (.A(_06267_),
    .Y(net4240));
 BUFx3_ASAP7_75t_R place4242 (.A(net4241),
    .Y(net4242));
 BUFx3_ASAP7_75t_R place4241 (.A(_06176_),
    .Y(net4241));
 BUFx3_ASAP7_75t_R place4243 (.A(_06149_),
    .Y(net4243));
 BUFx3_ASAP7_75t_R place4244 (.A(_06094_),
    .Y(net4244));
 BUFx3_ASAP7_75t_R place4245 (.A(_06048_),
    .Y(net4245));
 BUFx3_ASAP7_75t_R place4255 (.A(_05478_),
    .Y(net4255));
 BUFx3_ASAP7_75t_R place4247 (.A(_05977_),
    .Y(net4247));
 BUFx3_ASAP7_75t_R place4248 (.A(_05915_),
    .Y(net4248));
 BUFx3_ASAP7_75t_R place4249 (.A(_05658_),
    .Y(net4249));
 BUFx3_ASAP7_75t_R place4250 (.A(_05577_),
    .Y(net4250));
 BUFx3_ASAP7_75t_R place4251 (.A(_05547_),
    .Y(net4251));
 BUFx3_ASAP7_75t_R place4252 (.A(net5960),
    .Y(net4252));
 BUFx3_ASAP7_75t_R place4253 (.A(_05491_),
    .Y(net4253));
 BUFx3_ASAP7_75t_R place4254 (.A(_05478_),
    .Y(net4254));
 BUFx3_ASAP7_75t_R place4257 (.A(_05253_),
    .Y(net4257));
 BUFx3_ASAP7_75t_R place4256 (.A(_05335_),
    .Y(net4256));
 BUFx3_ASAP7_75t_R place4262 (.A(_05010_),
    .Y(net4262));
 BUFx3_ASAP7_75t_R place4263 (.A(_04724_),
    .Y(net4263));
 BUFx3_ASAP7_75t_R place4264 (.A(_04475_),
    .Y(net4264));
 BUFx3_ASAP7_75t_R place4265 (.A(_04469_),
    .Y(net4265));
 BUFx3_ASAP7_75t_R place4266 (.A(_04448_),
    .Y(net4266));
 BUFx3_ASAP7_75t_R place4276 (.A(net4275),
    .Y(net4276));
 BUFx3_ASAP7_75t_R place4267 (.A(_04409_),
    .Y(net4267));
 BUFx3_ASAP7_75t_R place4268 (.A(_04367_),
    .Y(net4268));
 BUFx3_ASAP7_75t_R place4269 (.A(_04288_),
    .Y(net4269));
 BUFx3_ASAP7_75t_R place4270 (.A(_03998_),
    .Y(net4270));
 BUFx3_ASAP7_75t_R place4271 (.A(_03920_),
    .Y(net4271));
 BUFx3_ASAP7_75t_R place4272 (.A(_03856_),
    .Y(net4272));
 BUFx3_ASAP7_75t_R place4273 (.A(_03600_),
    .Y(net4273));
 BUFx3_ASAP7_75t_R place4274 (.A(_03543_),
    .Y(net4274));
 BUFx3_ASAP7_75t_R place4275 (.A(_03289_),
    .Y(net4275));
 BUFx3_ASAP7_75t_R place4287 (.A(net4286),
    .Y(net4287));
 BUFx3_ASAP7_75t_R place4277 (.A(_03246_),
    .Y(net4277));
 BUFx3_ASAP7_75t_R place4285 (.A(_01330_),
    .Y(net4285));
 BUFx3_ASAP7_75t_R place4278 (.A(_03185_),
    .Y(net4278));
 BUFx3_ASAP7_75t_R place4279 (.A(_02762_),
    .Y(net4279));
 BUFx3_ASAP7_75t_R place4280 (.A(_02511_),
    .Y(net4280));
 BUFx3_ASAP7_75t_R place4281 (.A(_01573_),
    .Y(net4281));
 BUFx3_ASAP7_75t_R place4282 (.A(net5386),
    .Y(net4282));
 BUFx3_ASAP7_75t_R place4283 (.A(_01479_),
    .Y(net4283));
 BUFx3_ASAP7_75t_R place4284 (.A(net5380),
    .Y(net4284));
 BUFx6f_ASAP7_75t_R place4286 (.A(_01077_),
    .Y(net4286));
 BUFx3_ASAP7_75t_R place4307 (.A(net4306),
    .Y(net4307));
 BUFx3_ASAP7_75t_R place4297 (.A(net4296),
    .Y(net4297));
 BUFx3_ASAP7_75t_R place4294 (.A(_06372_),
    .Y(net4294));
 BUFx3_ASAP7_75t_R place4292 (.A(_06445_),
    .Y(net4292));
 BUFx3_ASAP7_75t_R place4291 (.A(_06464_),
    .Y(net4291));
 BUFx3_ASAP7_75t_R place4293 (.A(_06399_),
    .Y(net4293));
 BUFx3_ASAP7_75t_R place4295 (.A(_06343_),
    .Y(net4295));
 BUFx3_ASAP7_75t_R place4296 (.A(_06272_),
    .Y(net4296));
 BUFx3_ASAP7_75t_R place4301 (.A(_06110_),
    .Y(net4301));
 BUFx3_ASAP7_75t_R place4298 (.A(_06266_),
    .Y(net4298));
 BUFx3_ASAP7_75t_R place4299 (.A(_06157_),
    .Y(net4299));
 BUFx3_ASAP7_75t_R place4300 (.A(_06110_),
    .Y(net4300));
 BUFx3_ASAP7_75t_R place4306 (.A(_05503_),
    .Y(net4306));
 BUFx3_ASAP7_75t_R place4303 (.A(_05599_),
    .Y(net4303));
 BUFx3_ASAP7_75t_R place4302 (.A(_05600_),
    .Y(net4302));
 BUFx3_ASAP7_75t_R place4304 (.A(_05598_),
    .Y(net4304));
 BUFx3_ASAP7_75t_R place4305 (.A(_05523_),
    .Y(net4305));
 BUFx3_ASAP7_75t_R place4308 (.A(_05490_),
    .Y(net4308));
 BUFx3_ASAP7_75t_R place4309 (.A(_05477_),
    .Y(net4309));
 BUFx3_ASAP7_75t_R place4311 (.A(_05306_),
    .Y(net4311));
 BUFx3_ASAP7_75t_R place4312 (.A(_05252_),
    .Y(net4312));
 BUFx3_ASAP7_75t_R place4313 (.A(_05172_),
    .Y(net4313));
 BUFx3_ASAP7_75t_R place4314 (.A(_04517_),
    .Y(net4314));
 BUFx3_ASAP7_75t_R place4315 (.A(_04473_),
    .Y(net4315));
 BUFx3_ASAP7_75t_R place4316 (.A(_04450_),
    .Y(net4316));
 BUFx3_ASAP7_75t_R place4317 (.A(_04444_),
    .Y(net4317));
 BUFx3_ASAP7_75t_R place4318 (.A(_04433_),
    .Y(net4318));
 BUFx3_ASAP7_75t_R place4341 (.A(net4340),
    .Y(net4341));
 BUFx12f_ASAP7_75t_R place4330 (.A(net4329),
    .Y(net4330));
 BUFx3_ASAP7_75t_R place4319 (.A(_04428_),
    .Y(net4319));
 BUFx3_ASAP7_75t_R place4320 (.A(_04416_),
    .Y(net4320));
 BUFx3_ASAP7_75t_R place4321 (.A(_04397_),
    .Y(net4321));
 BUFx3_ASAP7_75t_R place4322 (.A(_04290_),
    .Y(net4322));
 BUFx6f_ASAP7_75t_R place4329 (.A(net4328),
    .Y(net4329));
 BUFx3_ASAP7_75t_R place4323 (.A(net5707),
    .Y(net4323));
 BUFx3_ASAP7_75t_R place4324 (.A(_03211_),
    .Y(net4324));
 BUFx3_ASAP7_75t_R place4325 (.A(_03201_),
    .Y(net4325));
 BUFx6f_ASAP7_75t_R place4326 (.A(_02761_),
    .Y(net4326));
 BUFx3_ASAP7_75t_R place4327 (.A(_02644_),
    .Y(net4327));
 BUFx6f_ASAP7_75t_R place4328 (.A(_02508_),
    .Y(net4328));
 BUFx3_ASAP7_75t_R place4331 (.A(_01575_),
    .Y(net4331));
 BUFx3_ASAP7_75t_R place4332 (.A(_01554_),
    .Y(net4332));
 BUFx3_ASAP7_75t_R place4333 (.A(_01467_),
    .Y(net4333));
 BUFx3_ASAP7_75t_R place4334 (.A(_01453_),
    .Y(net4334));
 BUFx3_ASAP7_75t_R place4335 (.A(net5918),
    .Y(net4335));
 BUFx3_ASAP7_75t_R place4336 (.A(net5428),
    .Y(net4336));
 BUFx3_ASAP7_75t_R place4337 (.A(_01412_),
    .Y(net4337));
 BUFx3_ASAP7_75t_R place4338 (.A(_01329_),
    .Y(net4338));
 BUFx3_ASAP7_75t_R place4339 (.A(_01281_),
    .Y(net4339));
 BUFx6f_ASAP7_75t_R place4340 (.A(_01076_),
    .Y(net4340));
 BUFx3_ASAP7_75t_R place4343 (.A(_05656_),
    .Y(net4343));
 BUFx3_ASAP7_75t_R place4344 (.A(_05616_),
    .Y(net4344));
 BUFx3_ASAP7_75t_R place4348 (.A(_05512_),
    .Y(net4348));
 BUFx3_ASAP7_75t_R place4345 (.A(_05576_),
    .Y(net4345));
 BUFx3_ASAP7_75t_R place4346 (.A(_05531_),
    .Y(net4346));
 BUFx3_ASAP7_75t_R place4347 (.A(_05515_),
    .Y(net4347));
 BUFx3_ASAP7_75t_R place4350 (.A(_04489_),
    .Y(net4350));
 BUFx3_ASAP7_75t_R place4351 (.A(_04480_),
    .Y(net4351));
 BUFx3_ASAP7_75t_R place4352 (.A(_04478_),
    .Y(net4352));
 BUFx3_ASAP7_75t_R place4354 (.A(_04454_),
    .Y(net4354));
 BUFx3_ASAP7_75t_R place4362 (.A(net4361),
    .Y(net4362));
 BUFx3_ASAP7_75t_R place4356 (.A(_04449_),
    .Y(net4356));
 BUFx3_ASAP7_75t_R place4357 (.A(_04442_),
    .Y(net4357));
 BUFx3_ASAP7_75t_R place4358 (.A(_04427_),
    .Y(net4358));
 BUFx3_ASAP7_75t_R place4359 (.A(_04415_),
    .Y(net4359));
 BUFx3_ASAP7_75t_R place4360 (.A(_04396_),
    .Y(net4360));
 BUFx6f_ASAP7_75t_R place4361 (.A(_04363_),
    .Y(net4361));
 BUFx3_ASAP7_75t_R place4369 (.A(_03203_),
    .Y(net4369));
 BUFx3_ASAP7_75t_R place4364 (.A(_04283_),
    .Y(net4364));
 BUFx3_ASAP7_75t_R place4365 (.A(_03267_),
    .Y(net4365));
 BUFx3_ASAP7_75t_R place4366 (.A(_03262_),
    .Y(net4366));
 BUFx3_ASAP7_75t_R place4367 (.A(_03254_),
    .Y(net4367));
 BUFx3_ASAP7_75t_R place4368 (.A(_03218_),
    .Y(net4368));
 BUFx3_ASAP7_75t_R place4370 (.A(_03200_),
    .Y(net4370));
 BUFx3_ASAP7_75t_R place4371 (.A(_02632_),
    .Y(net4371));
 BUFx3_ASAP7_75t_R place4372 (.A(_02507_),
    .Y(net4372));
 BUFx3_ASAP7_75t_R place4373 (.A(net5731),
    .Y(net4373));
 BUFx3_ASAP7_75t_R place4374 (.A(_00020_),
    .Y(net4374));
 BUFx3_ASAP7_75t_R place4375 (.A(_03038_),
    .Y(net4375));
 BUFx3_ASAP7_75t_R place4376 (.A(_01537_),
    .Y(net4376));
 BUFx3_ASAP7_75t_R place4377 (.A(_01534_),
    .Y(net4377));
 BUFx3_ASAP7_75t_R place4378 (.A(_01490_),
    .Y(net4378));
 BUFx3_ASAP7_75t_R place4379 (.A(_01475_),
    .Y(net4379));
 BUFx3_ASAP7_75t_R place4380 (.A(net5913),
    .Y(net4380));
 BUFx3_ASAP7_75t_R place4381 (.A(net5426),
    .Y(net4381));
 BUFx3_ASAP7_75t_R place4392 (.A(_05575_),
    .Y(net4392));
 BUFx3_ASAP7_75t_R place4382 (.A(_01445_),
    .Y(net4382));
 BUFx3_ASAP7_75t_R place4383 (.A(_01440_),
    .Y(net4383));
 BUFx3_ASAP7_75t_R place4384 (.A(net5385),
    .Y(net4384));
 BUFx3_ASAP7_75t_R place4385 (.A(_01415_),
    .Y(net4385));
 BUFx3_ASAP7_75t_R place4386 (.A(_01411_),
    .Y(net4386));
 BUFx3_ASAP7_75t_R place4387 (.A(_01408_),
    .Y(net4387));
 BUFx3_ASAP7_75t_R place4389 (.A(_01382_),
    .Y(net4389));
 BUFx3_ASAP7_75t_R place4388 (.A(_01387_),
    .Y(net4388));
 BUFx3_ASAP7_75t_R place4390 (.A(net5427),
    .Y(net4390));
 BUFx3_ASAP7_75t_R place4391 (.A(_05581_),
    .Y(net4391));
 BUFx3_ASAP7_75t_R place4393 (.A(_05564_),
    .Y(net4393));
 BUFx3_ASAP7_75t_R place4394 (.A(_05562_),
    .Y(net4394));
 BUFx3_ASAP7_75t_R place4395 (.A(_05535_),
    .Y(net4395));
 BUFx3_ASAP7_75t_R place4396 (.A(_05530_),
    .Y(net4396));
 BUFx3_ASAP7_75t_R place4398 (.A(_05514_),
    .Y(net4398));
 BUFx3_ASAP7_75t_R place4399 (.A(_05505_),
    .Y(net4399));
 BUFx12f_ASAP7_75t_R place4400 (.A(_05472_),
    .Y(net4400));
 BUFx3_ASAP7_75t_R place4424 (.A(_03253_),
    .Y(net4424));
 BUFx3_ASAP7_75t_R place4409 (.A(net4408),
    .Y(net4409));
 BUFx3_ASAP7_75t_R place4403 (.A(_04471_),
    .Y(net4403));
 BUFx3_ASAP7_75t_R place4404 (.A(_04452_),
    .Y(net4404));
 BUFx3_ASAP7_75t_R place4405 (.A(_04447_),
    .Y(net4405));
 BUFx3_ASAP7_75t_R place4406 (.A(_04445_),
    .Y(net4406));
 BUFx3_ASAP7_75t_R place4407 (.A(_04441_),
    .Y(net4407));
 BUFx3_ASAP7_75t_R place4408 (.A(_04426_),
    .Y(net4408));
 BUFx3_ASAP7_75t_R place4421 (.A(_03277_),
    .Y(net4421));
 BUFx3_ASAP7_75t_R place4410 (.A(_04412_),
    .Y(net4410));
 BUFx3_ASAP7_75t_R place4411 (.A(_04408_),
    .Y(net4411));
 BUFx3_ASAP7_75t_R place4412 (.A(_04403_),
    .Y(net4412));
 BUFx3_ASAP7_75t_R place4413 (.A(_04393_),
    .Y(net4413));
 BUFx3_ASAP7_75t_R place4414 (.A(_04384_),
    .Y(net4414));
 BUFx3_ASAP7_75t_R place4415 (.A(_04362_),
    .Y(net4415));
 BUFx3_ASAP7_75t_R place4416 (.A(_04361_),
    .Y(net4416));
 BUFx3_ASAP7_75t_R place4417 (.A(_04277_),
    .Y(net4417));
 BUFx3_ASAP7_75t_R place4418 (.A(_03317_),
    .Y(net4418));
 BUFx3_ASAP7_75t_R place4419 (.A(_03308_),
    .Y(net4419));
 BUFx3_ASAP7_75t_R place4420 (.A(_03281_),
    .Y(net4420));
 BUFx3_ASAP7_75t_R place4422 (.A(_03261_),
    .Y(net4422));
 BUFx3_ASAP7_75t_R place4423 (.A(_03257_),
    .Y(net4423));
 BUFx3_ASAP7_75t_R place4426 (.A(net5714),
    .Y(net4426));
 BUFx3_ASAP7_75t_R place4428 (.A(_03187_),
    .Y(net4428));
 BUFx3_ASAP7_75t_R place4429 (.A(_03134_),
    .Y(net4429));
 BUFx3_ASAP7_75t_R place4446 (.A(net4445),
    .Y(net4446));
 BUFx3_ASAP7_75t_R place4432 (.A(_01001_),
    .Y(net4432));
 BUFx3_ASAP7_75t_R place4442 (.A(_01335_),
    .Y(net4442));
 BUFx3_ASAP7_75t_R place4433 (.A(_01448_),
    .Y(net4433));
 BUFx3_ASAP7_75t_R place4434 (.A(_01426_),
    .Y(net4434));
 BUFx3_ASAP7_75t_R place4435 (.A(net5917),
    .Y(net4435));
 BUFx3_ASAP7_75t_R place4436 (.A(_01421_),
    .Y(net4436));
 BUFx3_ASAP7_75t_R place4437 (.A(_01420_),
    .Y(net4437));
 BUFx3_ASAP7_75t_R place4438 (.A(_01416_),
    .Y(net4438));
 BUFx3_ASAP7_75t_R place4439 (.A(_01407_),
    .Y(net4439));
 BUFx3_ASAP7_75t_R place4440 (.A(_01406_),
    .Y(net4440));
 BUFx3_ASAP7_75t_R place4441 (.A(_01383_),
    .Y(net4441));
 BUFx3_ASAP7_75t_R place4443 (.A(_01328_),
    .Y(net4443));
 BUFx3_ASAP7_75t_R place4444 (.A(_01322_),
    .Y(net4444));
 BUFx6f_ASAP7_75t_R place4445 (.A(_01260_),
    .Y(net4445));
 BUFx3_ASAP7_75t_R place4592 (.A(_01193_),
    .Y(net4592));
 BUFx3_ASAP7_75t_R place4447 (.A(_01247_),
    .Y(net4447));
 BUFx3_ASAP7_75t_R place4448 (.A(_01171_),
    .Y(net4448));
 BUFx3_ASAP7_75t_R place4460 (.A(net4459),
    .Y(net4460));
 BUFx3_ASAP7_75t_R place4450 (.A(_05519_),
    .Y(net4450));
 BUFx3_ASAP7_75t_R place4449 (.A(_05561_),
    .Y(net4449));
 BUFx3_ASAP7_75t_R place4451 (.A(_05509_),
    .Y(net4451));
 BUFx3_ASAP7_75t_R place4452 (.A(_05504_),
    .Y(net4452));
 BUFx3_ASAP7_75t_R place4456 (.A(net4455),
    .Y(net4456));
 BUFx3_ASAP7_75t_R place4453 (.A(_05489_),
    .Y(net4453));
 BUFx3_ASAP7_75t_R place4454 (.A(_05485_),
    .Y(net4454));
 BUFx3_ASAP7_75t_R place4455 (.A(_05471_),
    .Y(net4455));
 BUFx3_ASAP7_75t_R place4457 (.A(_04470_),
    .Y(net4457));
 BUFx6f_ASAP7_75t_R place4458 (.A(_04429_),
    .Y(net4458));
 BUFx6f_ASAP7_75t_R place4459 (.A(_04420_),
    .Y(net4459));
 BUFx6f_ASAP7_75t_R place4586 (.A(_01262_),
    .Y(net4586));
 BUFx3_ASAP7_75t_R place4464 (.A(_04246_),
    .Y(net4464));
 BUFx3_ASAP7_75t_R place4461 (.A(_04405_),
    .Y(net4461));
 BUFx3_ASAP7_75t_R place4462 (.A(_04402_),
    .Y(net4462));
 BUFx3_ASAP7_75t_R place4463 (.A(_04265_),
    .Y(net4463));
 BUFx3_ASAP7_75t_R place4585 (.A(_01262_),
    .Y(net4585));
 BUFx3_ASAP7_75t_R place4465 (.A(_03269_),
    .Y(net4465));
 BUFx3_ASAP7_75t_R place4466 (.A(_03259_),
    .Y(net4466));
 BUFx3_ASAP7_75t_R place4467 (.A(_03255_),
    .Y(net4467));
 BUFx3_ASAP7_75t_R place4468 (.A(_03244_),
    .Y(net4468));
 BUFx3_ASAP7_75t_R place4469 (.A(_03224_),
    .Y(net4469));
 BUFx3_ASAP7_75t_R place4581 (.A(_01360_),
    .Y(net4581));
 BUFx3_ASAP7_75t_R place4470 (.A(_03032_),
    .Y(net4470));
 BUFx3_ASAP7_75t_R place4471 (.A(_02557_),
    .Y(net4471));
 BUFx3_ASAP7_75t_R place4472 (.A(_02504_),
    .Y(net4472));
 BUFx3_ASAP7_75t_R place4575 (.A(_02706_),
    .Y(net4575));
 BUFx3_ASAP7_75t_R place4473 (.A(_03026_),
    .Y(net4473));
 BUFx3_ASAP7_75t_R place4474 (.A(_01424_),
    .Y(net4474));
 BUFx3_ASAP7_75t_R place4475 (.A(_01423_),
    .Y(net4475));
 BUFx3_ASAP7_75t_R place4476 (.A(_01419_),
    .Y(net4476));
 BUFx6f_ASAP7_75t_R place4570 (.A(_03059_),
    .Y(net4570));
 BUFx3_ASAP7_75t_R place4477 (.A(_01341_),
    .Y(net4477));
 BUFx3_ASAP7_75t_R place4478 (.A(net5379),
    .Y(net4478));
 BUFx3_ASAP7_75t_R place4479 (.A(_01327_),
    .Y(net4479));
 BUFx3_ASAP7_75t_R place4560 (.A(_03250_),
    .Y(net4560));
 BUFx3_ASAP7_75t_R place4480 (.A(_01316_),
    .Y(net4480));
 BUFx3_ASAP7_75t_R place4481 (.A(_01310_),
    .Y(net4481));
 BUFx3_ASAP7_75t_R place4528 (.A(_02598_),
    .Y(net4528));
 BUFx3_ASAP7_75t_R place4482 (.A(net5384),
    .Y(net4482));
 BUFx3_ASAP7_75t_R place4506 (.A(net4505),
    .Y(net4506));
 BUFx3_ASAP7_75t_R place4483 (.A(_01278_),
    .Y(net4483));
 BUFx3_ASAP7_75t_R place4484 (.A(_01274_),
    .Y(net4484));
 BUFx3_ASAP7_75t_R place4485 (.A(net5429),
    .Y(net4485));
 BUFx3_ASAP7_75t_R place4486 (.A(_01254_),
    .Y(net4486));
 BUFx3_ASAP7_75t_R place4487 (.A(_01253_),
    .Y(net4487));
 BUFx3_ASAP7_75t_R place4488 (.A(_01246_),
    .Y(net4488));
 BUFx3_ASAP7_75t_R place4489 (.A(_01245_),
    .Y(net4489));
 BUFx3_ASAP7_75t_R place4490 (.A(_01229_),
    .Y(net4490));
 BUFx3_ASAP7_75t_R place4491 (.A(_01228_),
    .Y(net4491));
 BUFx3_ASAP7_75t_R place4492 (.A(_01211_),
    .Y(net4492));
 BUFx3_ASAP7_75t_R place4493 (.A(_01210_),
    .Y(net4493));
 BUFx3_ASAP7_75t_R place4494 (.A(_01157_),
    .Y(net4494));
 BUFx3_ASAP7_75t_R place4502 (.A(_05484_),
    .Y(net4502));
 BUFx3_ASAP7_75t_R place4495 (.A(_05615_),
    .Y(net4495));
 BUFx3_ASAP7_75t_R place4496 (.A(_05582_),
    .Y(net4496));
 BUFx3_ASAP7_75t_R place4497 (.A(_05567_),
    .Y(net4497));
 BUFx3_ASAP7_75t_R place4499 (.A(net4498),
    .Y(net4499));
 BUFx6f_ASAP7_75t_R place4498 (.A(_05506_),
    .Y(net4498));
 BUFx3_ASAP7_75t_R place4500 (.A(_05499_),
    .Y(net4500));
 BUFx3_ASAP7_75t_R place4501 (.A(_05488_),
    .Y(net4501));
 BUFx3_ASAP7_75t_R place4503 (.A(_05479_),
    .Y(net4503));
 BUFx3_ASAP7_75t_R place4504 (.A(_05470_),
    .Y(net4504));
 BUFx3_ASAP7_75t_R place4505 (.A(_05469_),
    .Y(net4505));
 BUFx3_ASAP7_75t_R place4507 (.A(_05444_),
    .Y(net4507));
 BUFx3_ASAP7_75t_R place4508 (.A(_05430_),
    .Y(net4508));
 BUFx3_ASAP7_75t_R place4509 (.A(_04455_),
    .Y(net4509));
 BUFx3_ASAP7_75t_R place4510 (.A(_04414_),
    .Y(net4510));
 BUFx3_ASAP7_75t_R place4511 (.A(_04401_),
    .Y(net4511));
 BUFx3_ASAP7_75t_R place4512 (.A(_04395_),
    .Y(net4512));
 BUFx3_ASAP7_75t_R place4513 (.A(_04389_),
    .Y(net4513));
 BUFx3_ASAP7_75t_R place4514 (.A(_04387_),
    .Y(net4514));
 BUFx3_ASAP7_75t_R place4515 (.A(_04383_),
    .Y(net4515));
 BUFx3_ASAP7_75t_R place4516 (.A(_04375_),
    .Y(net4516));
 BUFx3_ASAP7_75t_R place4517 (.A(_04372_),
    .Y(net4517));
 BUFx3_ASAP7_75t_R place4518 (.A(_04356_),
    .Y(net4518));
 BUFx3_ASAP7_75t_R place4523 (.A(net4522),
    .Y(net4523));
 BUFx3_ASAP7_75t_R place4519 (.A(_03271_),
    .Y(net4519));
 BUFx3_ASAP7_75t_R place4520 (.A(_03256_),
    .Y(net4520));
 BUFx3_ASAP7_75t_R place4521 (.A(_03237_),
    .Y(net4521));
 BUFx3_ASAP7_75t_R place4522 (.A(_03223_),
    .Y(net4522));
 BUFx3_ASAP7_75t_R place4524 (.A(_03197_),
    .Y(net4524));
 BUFx3_ASAP7_75t_R place4525 (.A(_03127_),
    .Y(net4525));
 BUFx3_ASAP7_75t_R place4526 (.A(_02997_),
    .Y(net4526));
 BUFx3_ASAP7_75t_R place4527 (.A(_02937_),
    .Y(net4527));
 BUFx3_ASAP7_75t_R place4559 (.A(_04215_),
    .Y(net4559));
 BUFx3_ASAP7_75t_R place4529 (.A(_01391_),
    .Y(net4529));
 BUFx3_ASAP7_75t_R place4530 (.A(_01366_),
    .Y(net4530));
 BUFx3_ASAP7_75t_R place4531 (.A(_01326_),
    .Y(net4531));
 BUFx3_ASAP7_75t_R place4532 (.A(_01313_),
    .Y(net4532));
 BUFx3_ASAP7_75t_R place4533 (.A(_01309_),
    .Y(net4533));
 BUFx3_ASAP7_75t_R place4534 (.A(net5433),
    .Y(net4534));
 BUFx3_ASAP7_75t_R place4535 (.A(_01291_),
    .Y(net4535));
 BUFx3_ASAP7_75t_R place4536 (.A(_01290_),
    .Y(net4536));
 BUFx3_ASAP7_75t_R place4537 (.A(_01177_),
    .Y(net4537));
 BUFx3_ASAP7_75t_R place4538 (.A(_01169_),
    .Y(net4538));
 BUFx3_ASAP7_75t_R place4541 (.A(_05551_),
    .Y(net4541));
 BUFx3_ASAP7_75t_R place4539 (.A(_05565_),
    .Y(net4539));
 BUFx3_ASAP7_75t_R place4540 (.A(_05551_),
    .Y(net4540));
 BUFx3_ASAP7_75t_R place4542 (.A(_05533_),
    .Y(net4542));
 BUFx3_ASAP7_75t_R place4558 (.A(_04219_),
    .Y(net4558));
 BUFx3_ASAP7_75t_R place4543 (.A(_05529_),
    .Y(net4543));
 BUFx6f_ASAP7_75t_R place4544 (.A(_05526_),
    .Y(net4544));
 BUFx3_ASAP7_75t_R place4557 (.A(_04235_),
    .Y(net4557));
 BUFx3_ASAP7_75t_R place4545 (.A(net5665),
    .Y(net4545));
 BUFx3_ASAP7_75t_R place4546 (.A(_05494_),
    .Y(net4546));
 BUFx3_ASAP7_75t_R place4547 (.A(_05483_),
    .Y(net4547));
 BUFx3_ASAP7_75t_R place4548 (.A(_05439_),
    .Y(net4548));
 BUFx3_ASAP7_75t_R place4549 (.A(_04413_),
    .Y(net4549));
 BUFx3_ASAP7_75t_R place4550 (.A(_04398_),
    .Y(net4550));
 BUFx3_ASAP7_75t_R place4551 (.A(_04394_),
    .Y(net4551));
 BUFx3_ASAP7_75t_R place4552 (.A(_04382_),
    .Y(net4552));
 BUFx3_ASAP7_75t_R place4553 (.A(_04380_),
    .Y(net4553));
 BUFx3_ASAP7_75t_R place4554 (.A(_04355_),
    .Y(net4554));
 BUFx3_ASAP7_75t_R place4555 (.A(_04345_),
    .Y(net4555));
 BUFx3_ASAP7_75t_R place4556 (.A(_04249_),
    .Y(net4556));
 BUFx3_ASAP7_75t_R place4561 (.A(_03243_),
    .Y(net4561));
 BUFx3_ASAP7_75t_R place4562 (.A(_03227_),
    .Y(net4562));
 BUFx3_ASAP7_75t_R place4563 (.A(_03214_),
    .Y(net4563));
 BUFx3_ASAP7_75t_R place4564 (.A(_03196_),
    .Y(net4564));
 BUFx3_ASAP7_75t_R place4565 (.A(_03184_),
    .Y(net4565));
 BUFx3_ASAP7_75t_R place4566 (.A(_03181_),
    .Y(net4566));
 BUFx3_ASAP7_75t_R place4567 (.A(_03125_),
    .Y(net4567));
 BUFx3_ASAP7_75t_R place4568 (.A(_03120_),
    .Y(net4568));
 BUFx3_ASAP7_75t_R place4569 (.A(_03059_),
    .Y(net4569));
 BUFx3_ASAP7_75t_R place4573 (.A(_02741_),
    .Y(net4573));
 BUFx3_ASAP7_75t_R place4571 (.A(_03020_),
    .Y(net4571));
 BUFx3_ASAP7_75t_R place4572 (.A(_02984_),
    .Y(net4572));
 BUFx3_ASAP7_75t_R place4574 (.A(_02711_),
    .Y(net4574));
 BUFx3_ASAP7_75t_R place4576 (.A(_02539_),
    .Y(net4576));
 BUFx3_ASAP7_75t_R place4577 (.A(_00996_),
    .Y(net4577));
 BUFx3_ASAP7_75t_R place4580 (.A(_01374_),
    .Y(net4580));
 BUFx3_ASAP7_75t_R place4578 (.A(_03016_),
    .Y(net4578));
 BUFx3_ASAP7_75t_R place4579 (.A(_01431_),
    .Y(net4579));
 BUFx3_ASAP7_75t_R place4582 (.A(_01325_),
    .Y(net4582));
 BUFx3_ASAP7_75t_R place4583 (.A(_01287_),
    .Y(net4583));
 BUFx3_ASAP7_75t_R place4584 (.A(_01266_),
    .Y(net4584));
 BUFx3_ASAP7_75t_R place4587 (.A(_01255_),
    .Y(net4587));
 BUFx3_ASAP7_75t_R place4588 (.A(_01250_),
    .Y(net4588));
 BUFx3_ASAP7_75t_R place4589 (.A(_01239_),
    .Y(net4589));
 BUFx3_ASAP7_75t_R place4590 (.A(_01222_),
    .Y(net4590));
 BUFx3_ASAP7_75t_R place4591 (.A(_01219_),
    .Y(net4591));
 BUFx3_ASAP7_75t_R place4596 (.A(_01155_),
    .Y(net4596));
 BUFx6f_ASAP7_75t_R place4655 (.A(_01150_),
    .Y(net4655));
 BUFx3_ASAP7_75t_R place4597 (.A(_01152_),
    .Y(net4597));
 BUFx3_ASAP7_75t_R place4598 (.A(_01146_),
    .Y(net4598));
 BUFx3_ASAP7_75t_R place4599 (.A(_01062_),
    .Y(net4599));
 BUFx6f_ASAP7_75t_R place4635 (.A(_02841_),
    .Y(net4635));
 BUFx6f_ASAP7_75t_R place4634 (.A(_02841_),
    .Y(net4634));
 BUFx3_ASAP7_75t_R place4633 (.A(_02841_),
    .Y(net4633));
 BUFx3_ASAP7_75t_R place4600 (.A(_05558_),
    .Y(net4600));
 BUFx3_ASAP7_75t_R place4601 (.A(_05513_),
    .Y(net4601));
 BUFx3_ASAP7_75t_R place4602 (.A(_05508_),
    .Y(net4602));
 BUFx3_ASAP7_75t_R place4603 (.A(_05476_),
    .Y(net4603));
 BUFx3_ASAP7_75t_R place4632 (.A(_02841_),
    .Y(net4632));
 BUFx3_ASAP7_75t_R place4604 (.A(_05447_),
    .Y(net4604));
 BUFx3_ASAP7_75t_R place4605 (.A(_05443_),
    .Y(net4605));
 BUFx3_ASAP7_75t_R place4609 (.A(_04385_),
    .Y(net4609));
 BUFx3_ASAP7_75t_R place4606 (.A(_05435_),
    .Y(net4606));
 BUFx3_ASAP7_75t_R place4607 (.A(_05428_),
    .Y(net4607));
 BUFx3_ASAP7_75t_R place4608 (.A(_04437_),
    .Y(net4608));
 BUFx3_ASAP7_75t_R place4610 (.A(_04381_),
    .Y(net4610));
 BUFx3_ASAP7_75t_R place4611 (.A(_04376_),
    .Y(net4611));
 BUFx3_ASAP7_75t_R place4612 (.A(_04370_),
    .Y(net4612));
 BUFx3_ASAP7_75t_R place4631 (.A(_02841_),
    .Y(net4631));
 BUFx6f_ASAP7_75t_R place4630 (.A(_02841_),
    .Y(net4630));
 BUFx3_ASAP7_75t_R place4613 (.A(_04344_),
    .Y(net4613));
 BUFx3_ASAP7_75t_R place4614 (.A(_04341_),
    .Y(net4614));
 BUFx3_ASAP7_75t_R place4615 (.A(_04225_),
    .Y(net4615));
 BUFx3_ASAP7_75t_R place4616 (.A(_04217_),
    .Y(net4616));
 BUFx3_ASAP7_75t_R place4617 (.A(_04214_),
    .Y(net4617));
 BUFx3_ASAP7_75t_R place4618 (.A(_03275_),
    .Y(net4618));
 BUFx3_ASAP7_75t_R place4619 (.A(_03260_),
    .Y(net4619));
 BUFx3_ASAP7_75t_R place4620 (.A(_03236_),
    .Y(net4620));
 BUFx3_ASAP7_75t_R place4621 (.A(_03234_),
    .Y(net4621));
 BUFx3_ASAP7_75t_R place4622 (.A(_03228_),
    .Y(net4622));
 BUFx3_ASAP7_75t_R place4627 (.A(_03057_),
    .Y(net4627));
 BUFx3_ASAP7_75t_R place4623 (.A(_03213_),
    .Y(net4623));
 BUFx6f_ASAP7_75t_R place4626 (.A(_03057_),
    .Y(net4626));
 BUFx3_ASAP7_75t_R place4624 (.A(_03116_),
    .Y(net4624));
 BUFx6f_ASAP7_75t_R place4625 (.A(_03057_),
    .Y(net4625));
 BUFx3_ASAP7_75t_R place4628 (.A(_03000_),
    .Y(net4628));
 BUFx3_ASAP7_75t_R place4629 (.A(_02983_),
    .Y(net4629));
 BUFx3_ASAP7_75t_R place4649 (.A(_01343_),
    .Y(net4649));
 BUFx3_ASAP7_75t_R place4641 (.A(_00973_),
    .Y(net4641));
 BUFx6f_ASAP7_75t_R place4639 (.A(_02497_),
    .Y(net4639));
 BUFx3_ASAP7_75t_R place4637 (.A(_02550_),
    .Y(net4637));
 BUFx3_ASAP7_75t_R place4636 (.A(_02705_),
    .Y(net4636));
 BUFx6f_ASAP7_75t_R place4647 (.A(_01373_),
    .Y(net4647));
 BUFx3_ASAP7_75t_R place4638 (.A(_02536_),
    .Y(net4638));
 BUFx3_ASAP7_75t_R place4640 (.A(_00994_),
    .Y(net4640));
 BUFx3_ASAP7_75t_R place4642 (.A(_00927_),
    .Y(net4642));
 BUFx3_ASAP7_75t_R place4643 (.A(_00490_),
    .Y(net4643));
 BUFx3_ASAP7_75t_R place4646 (.A(_01377_),
    .Y(net4646));
 BUFx3_ASAP7_75t_R place4644 (.A(_00355_),
    .Y(net4644));
 BUFx3_ASAP7_75t_R place4645 (.A(_01389_),
    .Y(net4645));
 BUFx3_ASAP7_75t_R place4648 (.A(_01348_),
    .Y(net4648));
 BUFx3_ASAP7_75t_R place4651 (.A(_01192_),
    .Y(net4651));
 BUFx3_ASAP7_75t_R place4650 (.A(_01204_),
    .Y(net4650));
 BUFx3_ASAP7_75t_R place4653 (.A(net5381),
    .Y(net4653));
 BUFx3_ASAP7_75t_R place4652 (.A(_01182_),
    .Y(net4652));
 BUFx3_ASAP7_75t_R place4654 (.A(_01154_),
    .Y(net4654));
 BUFx3_ASAP7_75t_R place5033 (.A(_01000_),
    .Y(net5033));
 BUFx6f_ASAP7_75t_R place5032 (.A(net5028),
    .Y(net5032));
 BUFx3_ASAP7_75t_R place5027 (.A(net5024),
    .Y(net5027));
 BUFx3_ASAP7_75t_R place4657 (.A(_01048_),
    .Y(net4657));
 BUFx3_ASAP7_75t_R place4696 (.A(_01132_),
    .Y(net4696));
 BUFx6f_ASAP7_75t_R place4695 (.A(_01132_),
    .Y(net4695));
 BUFx3_ASAP7_75t_R place4694 (.A(net4693),
    .Y(net4694));
 BUFx6f_ASAP7_75t_R place4693 (.A(_01132_),
    .Y(net4693));
 BUFx3_ASAP7_75t_R place4674 (.A(_04212_),
    .Y(net4674));
 BUFx3_ASAP7_75t_R place4662 (.A(_05463_),
    .Y(net4662));
 BUFx3_ASAP7_75t_R place4658 (.A(_00464_),
    .Y(net4658));
 BUFx3_ASAP7_75t_R place4659 (.A(_00339_),
    .Y(net4659));
 BUFx3_ASAP7_75t_R place4660 (.A(_05507_),
    .Y(net4660));
 BUFx3_ASAP7_75t_R place4661 (.A(_05482_),
    .Y(net4661));
 BUFx3_ASAP7_75t_R place4663 (.A(_05442_),
    .Y(net4663));
 BUFx3_ASAP7_75t_R place4664 (.A(_05437_),
    .Y(net4664));
 BUFx3_ASAP7_75t_R place4665 (.A(_05434_),
    .Y(net4665));
 BUFx3_ASAP7_75t_R place4666 (.A(net5604),
    .Y(net4666));
 BUFx3_ASAP7_75t_R place4667 (.A(_04369_),
    .Y(net4667));
 BUFx3_ASAP7_75t_R place4668 (.A(_04366_),
    .Y(net4668));
 BUFx3_ASAP7_75t_R place4669 (.A(_04350_),
    .Y(net4669));
 BUFx3_ASAP7_75t_R place4670 (.A(_04343_),
    .Y(net4670));
 BUFx3_ASAP7_75t_R place4671 (.A(_04338_),
    .Y(net4671));
 BUFx3_ASAP7_75t_R place4672 (.A(_04213_),
    .Y(net4672));
 BUFx3_ASAP7_75t_R place4673 (.A(_04212_),
    .Y(net4673));
 BUFx3_ASAP7_75t_R place4683 (.A(_02977_),
    .Y(net4683));
 BUFx3_ASAP7_75t_R place4675 (.A(_03274_),
    .Y(net4675));
 BUFx3_ASAP7_75t_R place4676 (.A(_03233_),
    .Y(net4676));
 BUFx3_ASAP7_75t_R place4677 (.A(_03220_),
    .Y(net4677));
 BUFx3_ASAP7_75t_R place4678 (.A(_03194_),
    .Y(net4678));
 BUFx3_ASAP7_75t_R place4679 (.A(_03174_),
    .Y(net4679));
 BUFx3_ASAP7_75t_R place4680 (.A(_03168_),
    .Y(net4680));
 BUFx3_ASAP7_75t_R place4681 (.A(_03115_),
    .Y(net4681));
 BUFx3_ASAP7_75t_R place4682 (.A(_02977_),
    .Y(net4682));
 BUFx6f_ASAP7_75t_R place4689 (.A(_02520_),
    .Y(net4689));
 BUFx3_ASAP7_75t_R place4684 (.A(_02805_),
    .Y(net4684));
 BUFx3_ASAP7_75t_R place4685 (.A(_02786_),
    .Y(net4685));
 BUFx3_ASAP7_75t_R place4686 (.A(_02549_),
    .Y(net4686));
 BUFx3_ASAP7_75t_R place4687 (.A(_02534_),
    .Y(net4687));
 BUFx6f_ASAP7_75t_R place4688 (.A(_02520_),
    .Y(net4688));
 BUFx3_ASAP7_75t_R place4690 (.A(_02513_),
    .Y(net4690));
 BUFx3_ASAP7_75t_R place4691 (.A(_02496_),
    .Y(net4691));
 BUFx3_ASAP7_75t_R place4692 (.A(_01132_),
    .Y(net4692));
 BUFx6f_ASAP7_75t_R place5026 (.A(net5024),
    .Y(net5026));
 BUFx3_ASAP7_75t_R place4697 (.A(_00993_),
    .Y(net4697));
 BUFx3_ASAP7_75t_R place4698 (.A(_00982_),
    .Y(net4698));
 BUFx3_ASAP7_75t_R place4699 (.A(_00972_),
    .Y(net4699));
 BUFx3_ASAP7_75t_R place4700 (.A(_00885_),
    .Y(net4700));
 BUFx3_ASAP7_75t_R place4701 (.A(_00463_),
    .Y(net4701));
 BUFx6f_ASAP7_75t_R place5025 (.A(net5024),
    .Y(net5025));
 BUFx3_ASAP7_75t_R place5024 (.A(_01003_),
    .Y(net5024));
 BUFx3_ASAP7_75t_R place4708 (.A(_01388_),
    .Y(net4708));
 BUFx3_ASAP7_75t_R place4702 (.A(_03039_),
    .Y(net4702));
 BUFx3_ASAP7_75t_R place4703 (.A(_03033_),
    .Y(net4703));
 BUFx3_ASAP7_75t_R place4704 (.A(_03027_),
    .Y(net4704));
 BUFx3_ASAP7_75t_R place4705 (.A(_03021_),
    .Y(net4705));
 BUFx3_ASAP7_75t_R place4706 (.A(_01401_),
    .Y(net4706));
 BUFx3_ASAP7_75t_R place4707 (.A(_01394_),
    .Y(net4707));
 BUFx3_ASAP7_75t_R place4709 (.A(_01363_),
    .Y(net4709));
 BUFx3_ASAP7_75t_R place4710 (.A(_01358_),
    .Y(net4710));
 BUFx3_ASAP7_75t_R place5023 (.A(net5022),
    .Y(net5023));
 BUFx3_ASAP7_75t_R place5011 (.A(net5010),
    .Y(net5011));
 BUFx3_ASAP7_75t_R place5000 (.A(\u_fft.sched[47] ),
    .Y(net5000));
 BUFx3_ASAP7_75t_R place4998 (.A(\u_fft.sched[48] ),
    .Y(net4998));
 BUFx3_ASAP7_75t_R place4921 (.A(_02541_),
    .Y(net4921));
 BUFx3_ASAP7_75t_R place4920 (.A(_02566_),
    .Y(net4920));
 BUFx3_ASAP7_75t_R place4915 (.A(_02599_),
    .Y(net4915));
 BUFx3_ASAP7_75t_R place4904 (.A(_02714_),
    .Y(net4904));
 BUFx3_ASAP7_75t_R place4902 (.A(_02753_),
    .Y(net4902));
 BUFx3_ASAP7_75t_R place4901 (.A(_02827_),
    .Y(net4901));
 BUFx3_ASAP7_75t_R place4900 (.A(_02924_),
    .Y(net4900));
 BUFx3_ASAP7_75t_R place4711 (.A(_01144_),
    .Y(net4711));
 BUFx3_ASAP7_75t_R place4712 (.A(_01069_),
    .Y(net4712));
 BUFx3_ASAP7_75t_R place4713 (.A(_01067_),
    .Y(net4713));
 BUFx3_ASAP7_75t_R place4899 (.A(_02929_),
    .Y(net4899));
 BUFx3_ASAP7_75t_R place4716 (.A(_01049_),
    .Y(net4716));
 BUFx3_ASAP7_75t_R place4715 (.A(_01049_),
    .Y(net4715));
 BUFx3_ASAP7_75t_R place4714 (.A(_01052_),
    .Y(net4714));
 BUFx3_ASAP7_75t_R place4898 (.A(_02990_),
    .Y(net4898));
 BUFx3_ASAP7_75t_R place4891 (.A(_03100_),
    .Y(net4891));
 BUFx3_ASAP7_75t_R place4894 (.A(_03083_),
    .Y(net4894));
 BUFx3_ASAP7_75t_R place4890 (.A(_03105_),
    .Y(net4890));
 BUFx6f_ASAP7_75t_R place4888 (.A(_03165_),
    .Y(net4888));
 BUFx3_ASAP7_75t_R place4761 (.A(net4760),
    .Y(net4761));
 BUFx3_ASAP7_75t_R place4758 (.A(net4757),
    .Y(net4758));
 BUFx3_ASAP7_75t_R place4754 (.A(_00532_),
    .Y(net4754));
 BUFx3_ASAP7_75t_R place4751 (.A(_00911_),
    .Y(net4751));
 BUFx3_ASAP7_75t_R place4749 (.A(_00978_),
    .Y(net4749));
 BUFx3_ASAP7_75t_R place4747 (.A(_01126_),
    .Y(net4747));
 BUFx3_ASAP7_75t_R place4740 (.A(_02738_),
    .Y(net4740));
 BUFx3_ASAP7_75t_R place4739 (.A(_02776_),
    .Y(net4739));
 BUFx3_ASAP7_75t_R place4737 (.A(net4736),
    .Y(net4737));
 BUFx3_ASAP7_75t_R place4735 (.A(_02936_),
    .Y(net4735));
 BUFx3_ASAP7_75t_R place4727 (.A(_04211_),
    .Y(net4727));
 BUFx3_ASAP7_75t_R place4717 (.A(_01014_),
    .Y(net4717));
 BUFx3_ASAP7_75t_R place4724 (.A(_04339_),
    .Y(net4724));
 BUFx6f_ASAP7_75t_R place4719 (.A(_05445_),
    .Y(net4719));
 BUFx3_ASAP7_75t_R place4718 (.A(_05496_),
    .Y(net4718));
 BUFx3_ASAP7_75t_R place4720 (.A(_05436_),
    .Y(net4720));
 BUFx3_ASAP7_75t_R place4721 (.A(_05433_),
    .Y(net4721));
 BUFx3_ASAP7_75t_R place4722 (.A(_05424_),
    .Y(net4722));
 BUFx3_ASAP7_75t_R place4723 (.A(_04349_),
    .Y(net4723));
 BUFx3_ASAP7_75t_R place4725 (.A(_04252_),
    .Y(net4725));
 BUFx3_ASAP7_75t_R place4726 (.A(_04234_),
    .Y(net4726));
 BUFx3_ASAP7_75t_R place4728 (.A(_04207_),
    .Y(net4728));
 BUFx3_ASAP7_75t_R place4729 (.A(_03191_),
    .Y(net4729));
 BUFx3_ASAP7_75t_R place4730 (.A(_03179_),
    .Y(net4730));
 BUFx3_ASAP7_75t_R place4731 (.A(_03178_),
    .Y(net4731));
 BUFx3_ASAP7_75t_R place4732 (.A(_03176_),
    .Y(net4732));
 BUFx3_ASAP7_75t_R place4733 (.A(_03172_),
    .Y(net4733));
 BUFx3_ASAP7_75t_R place4734 (.A(_03096_),
    .Y(net4734));
 BUFx6f_ASAP7_75t_R place4736 (.A(_02894_),
    .Y(net4736));
 BUFx3_ASAP7_75t_R place4738 (.A(_02785_),
    .Y(net4738));
 BUFx3_ASAP7_75t_R place4741 (.A(_02735_),
    .Y(net4741));
 BUFx3_ASAP7_75t_R place4742 (.A(_02548_),
    .Y(net4742));
 BUFx3_ASAP7_75t_R place4743 (.A(_02533_),
    .Y(net4743));
 BUFx3_ASAP7_75t_R place4744 (.A(net5692),
    .Y(net4744));
 BUFx3_ASAP7_75t_R place4745 (.A(_00487_),
    .Y(net4745));
 BUFx3_ASAP7_75t_R place4746 (.A(_01131_),
    .Y(net4746));
 BUFx3_ASAP7_75t_R place4748 (.A(_00986_),
    .Y(net4748));
 BUFx3_ASAP7_75t_R place4750 (.A(_00951_),
    .Y(net4750));
 BUFx3_ASAP7_75t_R place4752 (.A(_00542_),
    .Y(net4752));
 BUFx3_ASAP7_75t_R place4753 (.A(_00540_),
    .Y(net4753));
 BUFx3_ASAP7_75t_R place4755 (.A(_00513_),
    .Y(net4755));
 BUFx3_ASAP7_75t_R place4756 (.A(_00503_),
    .Y(net4756));
 BUFx3_ASAP7_75t_R place4757 (.A(_00501_),
    .Y(net4757));
 BUFx3_ASAP7_75t_R place4760 (.A(_00462_),
    .Y(net4760));
 BUFx3_ASAP7_75t_R place4759 (.A(_00469_),
    .Y(net4759));
 BUFx3_ASAP7_75t_R place4884 (.A(_04222_),
    .Y(net4884));
 BUFx3_ASAP7_75t_R place4762 (.A(net5365),
    .Y(net4762));
 BUFx3_ASAP7_75t_R place4871 (.A(_05480_),
    .Y(net4871));
 BUFx3_ASAP7_75t_R place4764 (.A(net4763),
    .Y(net4764));
 BUFx3_ASAP7_75t_R place4763 (.A(_00456_),
    .Y(net4763));
 BUFx3_ASAP7_75t_R place4868 (.A(_00527_),
    .Y(net4868));
 BUFx3_ASAP7_75t_R place4801 (.A(net5366),
    .Y(net4801));
 BUFx3_ASAP7_75t_R place4765 (.A(_00454_),
    .Y(net4765));
 BUFx3_ASAP7_75t_R place4768 (.A(net5393),
    .Y(net4768));
 BUFx3_ASAP7_75t_R place4766 (.A(_00452_),
    .Y(net4766));
 BUFx3_ASAP7_75t_R place4767 (.A(_00450_),
    .Y(net4767));
 BUFx3_ASAP7_75t_R place4770 (.A(net4769),
    .Y(net4770));
 BUFx3_ASAP7_75t_R place4769 (.A(_00448_),
    .Y(net4769));
 BUFx3_ASAP7_75t_R place4772 (.A(net5436),
    .Y(net4772));
 BUFx3_ASAP7_75t_R place4771 (.A(_00446_),
    .Y(net4771));
 BUFx3_ASAP7_75t_R place4774 (.A(net4773),
    .Y(net4774));
 BUFx3_ASAP7_75t_R place4773 (.A(_00444_),
    .Y(net4773));
 BUFx3_ASAP7_75t_R place4776 (.A(net4775),
    .Y(net4776));
 BUFx3_ASAP7_75t_R place4775 (.A(_00442_),
    .Y(net4775));
 BUFx3_ASAP7_75t_R place4778 (.A(net4777),
    .Y(net4778));
 BUFx3_ASAP7_75t_R place4777 (.A(_00440_),
    .Y(net4777));
 BUFx3_ASAP7_75t_R place4780 (.A(net4779),
    .Y(net4780));
 BUFx6f_ASAP7_75t_R place4779 (.A(net5367),
    .Y(net4779));
 BUFx3_ASAP7_75t_R place4782 (.A(net4781),
    .Y(net4782));
 BUFx3_ASAP7_75t_R place4781 (.A(_00436_),
    .Y(net4781));
 BUFx3_ASAP7_75t_R place4784 (.A(net4783),
    .Y(net4784));
 BUFx3_ASAP7_75t_R place4783 (.A(_00434_),
    .Y(net4783));
 BUFx3_ASAP7_75t_R place4786 (.A(net4785),
    .Y(net4786));
 BUFx3_ASAP7_75t_R place4785 (.A(_00432_),
    .Y(net4785));
 BUFx3_ASAP7_75t_R place4788 (.A(net4787),
    .Y(net4788));
 BUFx3_ASAP7_75t_R place4787 (.A(_00430_),
    .Y(net4787));
 BUFx3_ASAP7_75t_R place4790 (.A(net4789),
    .Y(net4790));
 BUFx3_ASAP7_75t_R place4789 (.A(_00428_),
    .Y(net4789));
 BUFx3_ASAP7_75t_R place4792 (.A(net4791),
    .Y(net4792));
 BUFx3_ASAP7_75t_R place4791 (.A(_00426_),
    .Y(net4791));
 BUFx3_ASAP7_75t_R place4794 (.A(net4793),
    .Y(net4794));
 BUFx3_ASAP7_75t_R place4793 (.A(_00424_),
    .Y(net4793));
 BUFx3_ASAP7_75t_R place4796 (.A(net4795),
    .Y(net4796));
 BUFx3_ASAP7_75t_R place4795 (.A(_00422_),
    .Y(net4795));
 BUFx3_ASAP7_75t_R place4798 (.A(net4797),
    .Y(net4798));
 BUFx3_ASAP7_75t_R place4797 (.A(_00420_),
    .Y(net4797));
 BUFx3_ASAP7_75t_R place4800 (.A(net4799),
    .Y(net4800));
 BUFx3_ASAP7_75t_R place4799 (.A(_00418_),
    .Y(net4799));
 BUFx3_ASAP7_75t_R place4803 (.A(net4802),
    .Y(net4803));
 BUFx3_ASAP7_75t_R place4802 (.A(_00416_),
    .Y(net4802));
 BUFx3_ASAP7_75t_R place4805 (.A(net4804),
    .Y(net4805));
 BUFx3_ASAP7_75t_R place4804 (.A(_00414_),
    .Y(net4804));
 BUFx3_ASAP7_75t_R place4807 (.A(net4806),
    .Y(net4807));
 BUFx3_ASAP7_75t_R place4806 (.A(_00412_),
    .Y(net4806));
 BUFx3_ASAP7_75t_R place4865 (.A(_00877_),
    .Y(net4865));
 BUFx3_ASAP7_75t_R place4809 (.A(net4808),
    .Y(net4809));
 BUFx3_ASAP7_75t_R place4808 (.A(_00410_),
    .Y(net4808));
 BUFx3_ASAP7_75t_R place4811 (.A(net5376),
    .Y(net4811));
 BUFx3_ASAP7_75t_R place4810 (.A(net5376),
    .Y(net4810));
 BUFx3_ASAP7_75t_R place4864 (.A(_00883_),
    .Y(net4864));
 BUFx3_ASAP7_75t_R place4860 (.A(_00950_),
    .Y(net4860));
 BUFx3_ASAP7_75t_R place4812 (.A(_00406_),
    .Y(net4812));
 BUFx3_ASAP7_75t_R place4851 (.A(_02564_),
    .Y(net4851));
 BUFx3_ASAP7_75t_R place4813 (.A(_00404_),
    .Y(net4813));
 BUFx3_ASAP7_75t_R place4850 (.A(_02732_),
    .Y(net4850));
 BUFx3_ASAP7_75t_R place4848 (.A(_02815_),
    .Y(net4848));
 BUFx3_ASAP7_75t_R place4814 (.A(_00552_),
    .Y(net4814));
 BUFx3_ASAP7_75t_R place4815 (.A(net5603),
    .Y(net4815));
 BUFx3_ASAP7_75t_R place4816 (.A(_00539_),
    .Y(net4816));
 BUFx3_ASAP7_75t_R place4817 (.A(net5710),
    .Y(net4817));
 BUFx3_ASAP7_75t_R place4818 (.A(_00531_),
    .Y(net4818));
 BUFx3_ASAP7_75t_R place4819 (.A(_00522_),
    .Y(net4819));
 BUFx3_ASAP7_75t_R place4820 (.A(_00516_),
    .Y(net4820));
 BUFx3_ASAP7_75t_R place4821 (.A(_00514_),
    .Y(net4821));
 BUFx3_ASAP7_75t_R place4822 (.A(_00468_),
    .Y(net4822));
 BUFx3_ASAP7_75t_R place4823 (.A(_00460_),
    .Y(net4823));
 BUFx3_ASAP7_75t_R place4824 (.A(_00457_),
    .Y(net4824));
 BUFx3_ASAP7_75t_R place4826 (.A(net4825),
    .Y(net4826));
 BUFx6f_ASAP7_75t_R place4825 (.A(_00455_),
    .Y(net4825));
 BUFx3_ASAP7_75t_R place4846 (.A(_02907_),
    .Y(net4846));
 BUFx3_ASAP7_75t_R place4827 (.A(_00453_),
    .Y(net4827));
 BUFx3_ASAP7_75t_R place4828 (.A(_00451_),
    .Y(net4828));
 BUFx3_ASAP7_75t_R place4840 (.A(_04223_),
    .Y(net4840));
 BUFx3_ASAP7_75t_R place4839 (.A(_04251_),
    .Y(net4839));
 BUFx3_ASAP7_75t_R place4829 (.A(_00443_),
    .Y(net4829));
 BUFx3_ASAP7_75t_R place4830 (.A(_00439_),
    .Y(net4830));
 BUFx3_ASAP7_75t_R place4833 (.A(_00409_),
    .Y(net4833));
 BUFx3_ASAP7_75t_R place4831 (.A(_00427_),
    .Y(net4831));
 BUFx3_ASAP7_75t_R place4832 (.A(_00415_),
    .Y(net4832));
 BUFx3_ASAP7_75t_R place4835 (.A(_00403_),
    .Y(net4835));
 BUFx3_ASAP7_75t_R place4834 (.A(_00405_),
    .Y(net4834));
 BUFx3_ASAP7_75t_R place4836 (.A(_05495_),
    .Y(net4836));
 BUFx3_ASAP7_75t_R place4837 (.A(_04357_),
    .Y(net4837));
 BUFx3_ASAP7_75t_R place4838 (.A(_04336_),
    .Y(net4838));
 BUFx3_ASAP7_75t_R place4841 (.A(_03171_),
    .Y(net4841));
 BUFx3_ASAP7_75t_R place4842 (.A(_02993_),
    .Y(net4842));
 BUFx3_ASAP7_75t_R place4844 (.A(_02939_),
    .Y(net4844));
 BUFx3_ASAP7_75t_R place4843 (.A(_02939_),
    .Y(net4843));
 BUFx3_ASAP7_75t_R place4845 (.A(_02935_),
    .Y(net4845));
 BUFx3_ASAP7_75t_R place4847 (.A(_02901_),
    .Y(net4847));
 BUFx3_ASAP7_75t_R place4849 (.A(_02775_),
    .Y(net4849));
 BUFx3_ASAP7_75t_R place4852 (.A(_02547_),
    .Y(net4852));
 BUFx3_ASAP7_75t_R place4853 (.A(_01136_),
    .Y(net4853));
 BUFx3_ASAP7_75t_R place4858 (.A(_00984_),
    .Y(net4858));
 BUFx3_ASAP7_75t_R place4854 (.A(_01103_),
    .Y(net4854));
 BUFx3_ASAP7_75t_R place4855 (.A(_01004_),
    .Y(net4855));
 BUFx3_ASAP7_75t_R place4856 (.A(_00991_),
    .Y(net4856));
 BUFx3_ASAP7_75t_R place4857 (.A(_00988_),
    .Y(net4857));
 BUFx3_ASAP7_75t_R place4859 (.A(_00975_),
    .Y(net4859));
 BUFx3_ASAP7_75t_R place4861 (.A(_00945_),
    .Y(net4861));
 BUFx3_ASAP7_75t_R place4862 (.A(_00901_),
    .Y(net4862));
 BUFx3_ASAP7_75t_R place4863 (.A(_00898_),
    .Y(net4863));
 BUFx3_ASAP7_75t_R place4866 (.A(_06528_),
    .Y(net4866));
 BUFx3_ASAP7_75t_R place4867 (.A(_00536_),
    .Y(net4867));
 BUFx3_ASAP7_75t_R place4869 (.A(_00482_),
    .Y(net4869));
 BUFx3_ASAP7_75t_R place4870 (.A(_00367_),
    .Y(net4870));
 BUFx3_ASAP7_75t_R place4883 (.A(_04238_),
    .Y(net4883));
 BUFx3_ASAP7_75t_R place4872 (.A(_05464_),
    .Y(net4872));
 BUFx3_ASAP7_75t_R place4873 (.A(_05460_),
    .Y(net4873));
 BUFx3_ASAP7_75t_R place4874 (.A(_05459_),
    .Y(net4874));
 BUFx3_ASAP7_75t_R place4875 (.A(_05456_),
    .Y(net4875));
 BUFx3_ASAP7_75t_R place4876 (.A(_05454_),
    .Y(net4876));
 BUFx3_ASAP7_75t_R place4877 (.A(_05453_),
    .Y(net4877));
 BUFx3_ASAP7_75t_R place4878 (.A(_05451_),
    .Y(net4878));
 BUFx3_ASAP7_75t_R place4880 (.A(_04359_),
    .Y(net4880));
 BUFx3_ASAP7_75t_R place4879 (.A(_04390_),
    .Y(net4879));
 BUFx3_ASAP7_75t_R place4881 (.A(_04351_),
    .Y(net4881));
 BUFx3_ASAP7_75t_R place4882 (.A(_04347_),
    .Y(net4882));
 BUFx3_ASAP7_75t_R place4885 (.A(_03192_),
    .Y(net4885));
 BUFx3_ASAP7_75t_R place4886 (.A(_03189_),
    .Y(net4886));
 BUFx3_ASAP7_75t_R place4887 (.A(_03165_),
    .Y(net4887));
 BUFx3_ASAP7_75t_R place4889 (.A(_03141_),
    .Y(net4889));
 BUFx3_ASAP7_75t_R place4892 (.A(_03094_),
    .Y(net4892));
 BUFx3_ASAP7_75t_R place4893 (.A(_03089_),
    .Y(net4893));
 BUFx3_ASAP7_75t_R place4895 (.A(_03077_),
    .Y(net4895));
 BUFx3_ASAP7_75t_R place4896 (.A(_03053_),
    .Y(net4896));
 BUFx3_ASAP7_75t_R place4897 (.A(_02990_),
    .Y(net4897));
 BUFx3_ASAP7_75t_R place4903 (.A(_02734_),
    .Y(net4903));
 BUFx3_ASAP7_75t_R place4905 (.A(_02709_),
    .Y(net4905));
 BUFx3_ASAP7_75t_R place4906 (.A(_02669_),
    .Y(net4906));
 BUFx3_ASAP7_75t_R place4907 (.A(_02645_),
    .Y(net4907));
 BUFx3_ASAP7_75t_R place4908 (.A(_02640_),
    .Y(net4908));
 BUFx3_ASAP7_75t_R place4909 (.A(_02633_),
    .Y(net4909));
 BUFx3_ASAP7_75t_R place4910 (.A(_02628_),
    .Y(net4910));
 BUFx3_ASAP7_75t_R place4911 (.A(_02623_),
    .Y(net4911));
 BUFx3_ASAP7_75t_R place4912 (.A(_02618_),
    .Y(net4912));
 BUFx3_ASAP7_75t_R place4913 (.A(_02613_),
    .Y(net4913));
 BUFx3_ASAP7_75t_R place4914 (.A(_02608_),
    .Y(net4914));
 BUFx3_ASAP7_75t_R place4916 (.A(_02592_),
    .Y(net4916));
 BUFx3_ASAP7_75t_R place4917 (.A(_02587_),
    .Y(net4917));
 BUFx3_ASAP7_75t_R place4918 (.A(_02576_),
    .Y(net4918));
 BUFx3_ASAP7_75t_R place4919 (.A(_02571_),
    .Y(net4919));
 BUFx3_ASAP7_75t_R place4925 (.A(_02532_),
    .Y(net4925));
 BUFx3_ASAP7_75t_R place4922 (.A(_02538_),
    .Y(net4922));
 BUFx3_ASAP7_75t_R place4923 (.A(_02537_),
    .Y(net4923));
 BUFx3_ASAP7_75t_R place4924 (.A(_02535_),
    .Y(net4924));
 BUFx3_ASAP7_75t_R place4926 (.A(_02531_),
    .Y(net4926));
 BUFx3_ASAP7_75t_R place4927 (.A(\u_fft.sched[56] ),
    .Y(net4927));
 BUFx3_ASAP7_75t_R place4928 (.A(\u_fft.sched[58] ),
    .Y(net4928));
 BUFx3_ASAP7_75t_R place4929 (.A(\u_fft.sched[59] ),
    .Y(net4929));
 BUFx3_ASAP7_75t_R place4930 (.A(\u_fft.sched[60] ),
    .Y(net4930));
 BUFx3_ASAP7_75t_R place4931 (.A(\u_fft.sched[61] ),
    .Y(net4931));
 BUFx3_ASAP7_75t_R place4997 (.A(\u_fft.sched[51] ),
    .Y(net4997));
 BUFx3_ASAP7_75t_R place4932 (.A(\u_fft.sched[63] ),
    .Y(net4932));
 BUFx6f_ASAP7_75t_R place4935 (.A(\u_window_buffer.read_ptr[1] ),
    .Y(net4935));
 BUFx3_ASAP7_75t_R place4933 (.A(_02518_),
    .Y(net4933));
 BUFx3_ASAP7_75t_R place4934 (.A(_02517_),
    .Y(net4934));
 BUFx3_ASAP7_75t_R place4936 (.A(\u_window_buffer.read_ptr[2] ),
    .Y(net4936));
 BUFx3_ASAP7_75t_R place4937 (.A(\u_window_buffer.read_ptr[3] ),
    .Y(net4937));
 BUFx3_ASAP7_75t_R place4938 (.A(\u_window_buffer.read_ptr[4] ),
    .Y(net4938));
 BUFx3_ASAP7_75t_R place4939 (.A(\u_window_buffer.read_ptr[5] ),
    .Y(net4939));
 BUFx3_ASAP7_75t_R place4940 (.A(net5457),
    .Y(net4940));
 BUFx3_ASAP7_75t_R place4941 (.A(\u_window_buffer.read_ptr[7] ),
    .Y(net4941));
 BUFx3_ASAP7_75t_R place4942 (.A(\u_window_buffer.read_ptr[8] ),
    .Y(net4942));
 BUFx3_ASAP7_75t_R place4943 (.A(\u_window_buffer.read_ptr[9] ),
    .Y(net4943));
 BUFx3_ASAP7_75t_R place4944 (.A(\u_window_buffer.read_ptr[10] ),
    .Y(net4944));
 BUFx3_ASAP7_75t_R place4945 (.A(\u_window_buffer.read_ptr[11] ),
    .Y(net4945));
 BUFx3_ASAP7_75t_R place4946 (.A(\u_window_buffer.read_ptr[12] ),
    .Y(net4946));
 BUFx3_ASAP7_75t_R place4947 (.A(\u_window_buffer.read_ptr[13] ),
    .Y(net4947));
 BUFx3_ASAP7_75t_R place4948 (.A(\u_window_buffer.read_ptr[15] ),
    .Y(net4948));
 BUFx3_ASAP7_75t_R place4949 (.A(\u_window_buffer.read_ptr[16] ),
    .Y(net4949));
 BUFx3_ASAP7_75t_R place4950 (.A(\u_window_buffer.read_ptr[17] ),
    .Y(net4950));
 BUFx3_ASAP7_75t_R place4951 (.A(\u_window_buffer.read_ptr[18] ),
    .Y(net4951));
 BUFx3_ASAP7_75t_R place4952 (.A(\u_window_buffer.read_ptr[19] ),
    .Y(net4952));
 BUFx3_ASAP7_75t_R place4953 (.A(\u_window_buffer.read_ptr[20] ),
    .Y(net4953));
 BUFx3_ASAP7_75t_R place4954 (.A(\u_window_buffer.read_ptr[21] ),
    .Y(net4954));
 BUFx3_ASAP7_75t_R place4955 (.A(\u_window_buffer.read_ptr[22] ),
    .Y(net4955));
 BUFx3_ASAP7_75t_R place4956 (.A(\u_window_buffer.read_ptr[23] ),
    .Y(net4956));
 BUFx3_ASAP7_75t_R place4957 (.A(\u_window_buffer.read_ptr[24] ),
    .Y(net4957));
 BUFx3_ASAP7_75t_R place4958 (.A(\u_window_buffer.read_ptr[25] ),
    .Y(net4958));
 BUFx3_ASAP7_75t_R place4959 (.A(\u_window_buffer.read_ptr[26] ),
    .Y(net4959));
 BUFx3_ASAP7_75t_R place4960 (.A(\u_window_buffer.read_ptr[27] ),
    .Y(net4960));
 BUFx3_ASAP7_75t_R place4961 (.A(\u_window_buffer.read_ptr[28] ),
    .Y(net4961));
 BUFx3_ASAP7_75t_R place4962 (.A(\u_window_buffer.read_ptr[29] ),
    .Y(net4962));
 BUFx3_ASAP7_75t_R place4963 (.A(\u_window_buffer.read_ptr[30] ),
    .Y(net4963));
 BUFx3_ASAP7_75t_R place4964 (.A(\u_window_buffer.internal_read_ptr[6] ),
    .Y(net4964));
 BUFx6f_ASAP7_75t_R place4965 (.A(\u_window_buffer.internal_read_ptr[5] ),
    .Y(net4965));
 BUFx3_ASAP7_75t_R place4966 (.A(\u_window_buffer.internal_read_ptr[4] ),
    .Y(net4966));
 BUFx3_ASAP7_75t_R place4967 (.A(\u_window_buffer.internal_read_ptr[3] ),
    .Y(net4967));
 BUFx3_ASAP7_75t_R place4968 (.A(net5914),
    .Y(net4968));
 BUFx3_ASAP7_75t_R place4969 (.A(_02493_),
    .Y(net4969));
 BUFx3_ASAP7_75t_R place4970 (.A(\u_window_buffer.internal_read_ptr[1] ),
    .Y(net4970));
 BUFx3_ASAP7_75t_R place4971 (.A(\u_window_buffer.internal_read_ptr[7] ),
    .Y(net4971));
 BUFx3_ASAP7_75t_R place4972 (.A(\u_window_buffer.internal_read_ptr[8] ),
    .Y(net4972));
 BUFx3_ASAP7_75t_R place4973 (.A(\u_window_buffer.internal_read_ptr[9] ),
    .Y(net4973));
 BUFx3_ASAP7_75t_R place4974 (.A(\u_window_buffer.internal_read_ptr[10] ),
    .Y(net4974));
 BUFx3_ASAP7_75t_R place4975 (.A(\u_window_buffer.internal_read_ptr[11] ),
    .Y(net4975));
 BUFx3_ASAP7_75t_R place4976 (.A(\u_window_buffer.internal_read_ptr[12] ),
    .Y(net4976));
 BUFx3_ASAP7_75t_R place4977 (.A(\u_window_buffer.internal_read_ptr[13] ),
    .Y(net4977));
 BUFx3_ASAP7_75t_R place4978 (.A(\u_window_buffer.internal_read_ptr[14] ),
    .Y(net4978));
 BUFx3_ASAP7_75t_R place4979 (.A(\u_window_buffer.internal_read_ptr[15] ),
    .Y(net4979));
 BUFx3_ASAP7_75t_R place4980 (.A(\u_window_buffer.internal_read_ptr[16] ),
    .Y(net4980));
 BUFx3_ASAP7_75t_R place4981 (.A(\u_window_buffer.internal_read_ptr[17] ),
    .Y(net4981));
 BUFx3_ASAP7_75t_R place4982 (.A(\u_window_buffer.internal_read_ptr[18] ),
    .Y(net4982));
 BUFx3_ASAP7_75t_R place4983 (.A(\u_window_buffer.internal_read_ptr[19] ),
    .Y(net4983));
 BUFx3_ASAP7_75t_R place4984 (.A(\u_window_buffer.internal_read_ptr[20] ),
    .Y(net4984));
 BUFx3_ASAP7_75t_R place4985 (.A(\u_window_buffer.internal_read_ptr[21] ),
    .Y(net4985));
 BUFx3_ASAP7_75t_R place4986 (.A(\u_window_buffer.internal_read_ptr[22] ),
    .Y(net4986));
 BUFx3_ASAP7_75t_R place4987 (.A(\u_window_buffer.internal_read_ptr[23] ),
    .Y(net4987));
 BUFx3_ASAP7_75t_R place4988 (.A(\u_window_buffer.internal_read_ptr[24] ),
    .Y(net4988));
 BUFx3_ASAP7_75t_R place4989 (.A(\u_window_buffer.internal_read_ptr[25] ),
    .Y(net4989));
 BUFx3_ASAP7_75t_R place4990 (.A(\u_window_buffer.internal_read_ptr[26] ),
    .Y(net4990));
 BUFx3_ASAP7_75t_R place4991 (.A(\u_window_buffer.internal_read_ptr[27] ),
    .Y(net4991));
 BUFx3_ASAP7_75t_R place4992 (.A(\u_window_buffer.internal_read_ptr[28] ),
    .Y(net4992));
 BUFx3_ASAP7_75t_R place4993 (.A(\u_window_buffer.internal_read_ptr[29] ),
    .Y(net4993));
 BUFx3_ASAP7_75t_R place4994 (.A(\u_window_buffer.internal_read_ptr[30] ),
    .Y(net4994));
 BUFx3_ASAP7_75t_R place4995 (.A(\u_hamming_window.frame_ptr[0] ),
    .Y(net4995));
 BUFx3_ASAP7_75t_R place4996 (.A(\u_fft.sched[52] ),
    .Y(net4996));
 BUFx3_ASAP7_75t_R place4999 (.A(\u_fft.sched[46] ),
    .Y(net4999));
 BUFx3_ASAP7_75t_R place5001 (.A(\u_dct.n_ptr[1] ),
    .Y(net5001));
 BUFx3_ASAP7_75t_R place5002 (.A(\u_dct.n_ptr[0] ),
    .Y(net5002));
 BUFx3_ASAP7_75t_R place5003 (.A(_02487_),
    .Y(net5003));
 BUFx3_ASAP7_75t_R place5004 (.A(_02477_),
    .Y(net5004));
 BUFx3_ASAP7_75t_R place5005 (.A(_02469_),
    .Y(net5005));
 BUFx3_ASAP7_75t_R place5006 (.A(_02463_),
    .Y(net5006));
 BUFx3_ASAP7_75t_R place5007 (.A(_02458_),
    .Y(net5007));
 BUFx3_ASAP7_75t_R place5008 (.A(_02454_),
    .Y(net5008));
 BUFx3_ASAP7_75t_R place5009 (.A(_02449_),
    .Y(net5009));
 BUFx3_ASAP7_75t_R place5010 (.A(_02445_),
    .Y(net5010));
 BUFx3_ASAP7_75t_R place5012 (.A(_02426_),
    .Y(net5012));
 BUFx3_ASAP7_75t_R place5013 (.A(_02407_),
    .Y(net5013));
 BUFx3_ASAP7_75t_R place5014 (.A(_02392_),
    .Y(net5014));
 BUFx3_ASAP7_75t_R place5015 (.A(_02389_),
    .Y(net5015));
 BUFx3_ASAP7_75t_R place5016 (.A(_01135_),
    .Y(net5016));
 BUFx3_ASAP7_75t_R place5017 (.A(_01123_),
    .Y(net5017));
 BUFx3_ASAP7_75t_R place5018 (.A(_01104_),
    .Y(net5018));
 BUFx3_ASAP7_75t_R place5019 (.A(\u_window_buffer.read_ptr[0] ),
    .Y(net5019));
 BUFx3_ASAP7_75t_R place5020 (.A(net5623),
    .Y(net5020));
 BUFx3_ASAP7_75t_R place5021 (.A(\u_window_buffer.write_ptr[0] ),
    .Y(net5021));
 BUFx3_ASAP7_75t_R place5022 (.A(_01003_),
    .Y(net5022));
 BUFx3_ASAP7_75t_R place5031 (.A(net5028),
    .Y(net5031));
 BUFx3_ASAP7_75t_R place5030 (.A(net5028),
    .Y(net5030));
 BUFx3_ASAP7_75t_R place5029 (.A(net5028),
    .Y(net5029));
 BUFx6f_ASAP7_75t_R place5028 (.A(_01000_),
    .Y(net5028));
 BUFx3_ASAP7_75t_R place5044 (.A(\u_hamming_window.frame_ptr[1] ),
    .Y(net5044));
 BUFx3_ASAP7_75t_R place5040 (.A(\tx_fifo.write_ptr[0] ),
    .Y(net5040));
 BUFx3_ASAP7_75t_R place5035 (.A(_00985_),
    .Y(net5035));
 BUFx3_ASAP7_75t_R place5034 (.A(_00987_),
    .Y(net5034));
 BUFx3_ASAP7_75t_R place5036 (.A(_00964_),
    .Y(net5036));
 BUFx3_ASAP7_75t_R place5037 (.A(_00962_),
    .Y(net5037));
 BUFx3_ASAP7_75t_R place5038 (.A(_00960_),
    .Y(net5038));
 BUFx3_ASAP7_75t_R place5039 (.A(\tx_fifo.write_ptr[1] ),
    .Y(net5039));
 BUFx3_ASAP7_75t_R place5041 (.A(_00956_),
    .Y(net5041));
 BUFx3_ASAP7_75t_R place5043 (.A(_00949_),
    .Y(net5043));
 BUFx3_ASAP7_75t_R place5042 (.A(_00955_),
    .Y(net5042));
 BUFx3_ASAP7_75t_R place5045 (.A(_00942_),
    .Y(net5045));
 BUFx3_ASAP7_75t_R place5046 (.A(_00938_),
    .Y(net5046));
 BUFx3_ASAP7_75t_R place5047 (.A(_00937_),
    .Y(net5047));
 BUFx3_ASAP7_75t_R place5048 (.A(_00930_),
    .Y(net5048));
 BUFx3_ASAP7_75t_R place5056 (.A(_00924_),
    .Y(net5056));
 BUFx3_ASAP7_75t_R place5057 (.A(_00922_),
    .Y(net5057));
 BUFx3_ASAP7_75t_R place5058 (.A(_00910_),
    .Y(net5058));
 BUFx3_ASAP7_75t_R place5061 (.A(_00906_),
    .Y(net5061));
 BUFx3_ASAP7_75t_R place5064 (.A(_00895_),
    .Y(net5064));
 BUFx3_ASAP7_75t_R place5065 (.A(_00894_),
    .Y(net5065));
 BUFx3_ASAP7_75t_R place5066 (.A(\u_fft.sched[40] ),
    .Y(net5066));
 BUFx3_ASAP7_75t_R place5067 (.A(\u_fft.sched[41] ),
    .Y(net5067));
 BUFx3_ASAP7_75t_R place5068 (.A(\u_fft.sched[42] ),
    .Y(net5068));
 BUFx3_ASAP7_75t_R place5083 (.A(_00030_),
    .Y(net5083));
 BUFx3_ASAP7_75t_R place5070 (.A(\u_fft.sched[30] ),
    .Y(net5070));
 BUFx3_ASAP7_75t_R place5071 (.A(\u_fft.sched[31] ),
    .Y(net5071));
 BUFx3_ASAP7_75t_R place5072 (.A(\u_fft.sched[32] ),
    .Y(net5072));
 BUFx3_ASAP7_75t_R place5073 (.A(\u_fft.sched[33] ),
    .Y(net5073));
 BUFx3_ASAP7_75t_R place5074 (.A(\u_fft.sched[34] ),
    .Y(net5074));
 BUFx3_ASAP7_75t_R place5075 (.A(\u_fft.sched[35] ),
    .Y(net5075));
 BUFx3_ASAP7_75t_R place5076 (.A(\u_fft.sched[36] ),
    .Y(net5076));
 BUFx3_ASAP7_75t_R place5077 (.A(\u_fft.sched[37] ),
    .Y(net5077));
 BUFx3_ASAP7_75t_R place5078 (.A(\u_fft.sched[38] ),
    .Y(net5078));
 BUFx3_ASAP7_75t_R place5082 (.A(_06527_),
    .Y(net5082));
 BUFx3_ASAP7_75t_R place5079 (.A(_00882_),
    .Y(net5079));
 BUFx3_ASAP7_75t_R place5080 (.A(_00876_),
    .Y(net5080));
 BUFx3_ASAP7_75t_R place5081 (.A(_00875_),
    .Y(net5081));
 BUFx3_ASAP7_75t_R place5084 (.A(_00029_),
    .Y(net5084));
 BUFx3_ASAP7_75t_R place5085 (.A(_00028_),
    .Y(net5085));
 BUFx3_ASAP7_75t_R place5086 (.A(_00027_),
    .Y(net5086));
 BUFx3_ASAP7_75t_R place5087 (.A(_00025_),
    .Y(net5087));
 BUFx3_ASAP7_75t_R place5093 (.A(_00060_),
    .Y(net5093));
 BUFx3_ASAP7_75t_R place5089 (.A(_00070_),
    .Y(net5089));
 BUFx3_ASAP7_75t_R place5090 (.A(_00053_),
    .Y(net5090));
 BUFx3_ASAP7_75t_R place5091 (.A(_00052_),
    .Y(net5091));
 BUFx3_ASAP7_75t_R place5092 (.A(_00060_),
    .Y(net5092));
 BUFx3_ASAP7_75t_R place5190 (.A(_00151_),
    .Y(net5190));
 BUFx3_ASAP7_75t_R place5094 (.A(_00051_),
    .Y(net5094));
 BUFx3_ASAP7_75t_R place5098 (.A(net5097),
    .Y(net5098));
 BUFx3_ASAP7_75t_R place5095 (.A(_00049_),
    .Y(net5095));
 BUFx3_ASAP7_75t_R place5096 (.A(_00048_),
    .Y(net5096));
 BUFx3_ASAP7_75t_R place5097 (.A(_00047_),
    .Y(net5097));
 BUFx3_ASAP7_75t_R place5099 (.A(_00045_),
    .Y(net5099));
 BUFx3_ASAP7_75t_R place5100 (.A(_00044_),
    .Y(net5100));
 BUFx3_ASAP7_75t_R place5111 (.A(_00034_),
    .Y(net5111));
 BUFx3_ASAP7_75t_R place5101 (.A(_00043_),
    .Y(net5101));
 BUFx3_ASAP7_75t_R place5102 (.A(_00042_),
    .Y(net5102));
 BUFx3_ASAP7_75t_R place5103 (.A(_00041_),
    .Y(net5103));
 BUFx3_ASAP7_75t_R place5104 (.A(_00071_),
    .Y(net5104));
 BUFx3_ASAP7_75t_R place5105 (.A(_00040_),
    .Y(net5105));
 BUFx3_ASAP7_75t_R place5106 (.A(_00039_),
    .Y(net5106));
 BUFx3_ASAP7_75t_R place5107 (.A(_00038_),
    .Y(net5107));
 BUFx3_ASAP7_75t_R place5108 (.A(_00037_),
    .Y(net5108));
 BUFx3_ASAP7_75t_R place5109 (.A(_00036_),
    .Y(net5109));
 BUFx3_ASAP7_75t_R place5110 (.A(_00035_),
    .Y(net5110));
 BUFx3_ASAP7_75t_R place5112 (.A(_00033_),
    .Y(net5112));
 BUFx3_ASAP7_75t_R place5113 (.A(_00032_),
    .Y(net5113));
 BUFx3_ASAP7_75t_R place5114 (.A(_00031_),
    .Y(net5114));
 BUFx3_ASAP7_75t_R place5115 (.A(_00872_),
    .Y(net5115));
 BUFx3_ASAP7_75t_R place5116 (.A(_00072_),
    .Y(net5116));
 BUFx3_ASAP7_75t_R place5117 (.A(_00073_),
    .Y(net5117));
 BUFx3_ASAP7_75t_R place5118 (.A(_00074_),
    .Y(net5118));
 BUFx3_ASAP7_75t_R place5119 (.A(_00075_),
    .Y(net5119));
 BUFx3_ASAP7_75t_R place5120 (.A(net5395),
    .Y(net5120));
 BUFx3_ASAP7_75t_R place5121 (.A(_00077_),
    .Y(net5121));
 BUFx3_ASAP7_75t_R place5122 (.A(net5761),
    .Y(net5122));
 BUFx3_ASAP7_75t_R place5123 (.A(_00080_),
    .Y(net5123));
 BUFx3_ASAP7_75t_R place5124 (.A(_00082_),
    .Y(net5124));
 BUFx3_ASAP7_75t_R place5125 (.A(_00084_),
    .Y(net5125));
 BUFx3_ASAP7_75t_R place5126 (.A(_00085_),
    .Y(net5126));
 BUFx3_ASAP7_75t_R place5127 (.A(_00088_),
    .Y(net5127));
 BUFx3_ASAP7_75t_R place5128 (.A(_00089_),
    .Y(net5128));
 BUFx3_ASAP7_75t_R place5129 (.A(_00090_),
    .Y(net5129));
 BUFx3_ASAP7_75t_R place5130 (.A(_00091_),
    .Y(net5130));
 BUFx3_ASAP7_75t_R place5131 (.A(_00092_),
    .Y(net5131));
 BUFx3_ASAP7_75t_R place5132 (.A(_00093_),
    .Y(net5132));
 BUFx3_ASAP7_75t_R place5133 (.A(_00094_),
    .Y(net5133));
 BUFx3_ASAP7_75t_R place5134 (.A(_00095_),
    .Y(net5134));
 BUFx3_ASAP7_75t_R place5135 (.A(_00096_),
    .Y(net5135));
 BUFx3_ASAP7_75t_R place5136 (.A(_00097_),
    .Y(net5136));
 BUFx3_ASAP7_75t_R place5137 (.A(_00098_),
    .Y(net5137));
 BUFx3_ASAP7_75t_R place5138 (.A(_00099_),
    .Y(net5138));
 BUFx3_ASAP7_75t_R place5139 (.A(net5585),
    .Y(net5139));
 BUFx3_ASAP7_75t_R place5140 (.A(_00101_),
    .Y(net5140));
 BUFx3_ASAP7_75t_R place5141 (.A(_00102_),
    .Y(net5141));
 BUFx3_ASAP7_75t_R place5142 (.A(_00103_),
    .Y(net5142));
 BUFx3_ASAP7_75t_R place5143 (.A(_00461_),
    .Y(net5143));
 BUFx3_ASAP7_75t_R place5144 (.A(_00104_),
    .Y(net5144));
 BUFx3_ASAP7_75t_R place5145 (.A(_00337_),
    .Y(net5145));
 BUFx3_ASAP7_75t_R place5146 (.A(_00105_),
    .Y(net5146));
 BUFx3_ASAP7_75t_R place5147 (.A(_00106_),
    .Y(net5147));
 BUFx3_ASAP7_75t_R place5148 (.A(_00107_),
    .Y(net5148));
 BUFx3_ASAP7_75t_R place5149 (.A(_00108_),
    .Y(net5149));
 BUFx3_ASAP7_75t_R place5150 (.A(_00109_),
    .Y(net5150));
 BUFx3_ASAP7_75t_R place5151 (.A(_00110_),
    .Y(net5151));
 BUFx3_ASAP7_75t_R place5173 (.A(_00136_),
    .Y(net5173));
 BUFx3_ASAP7_75t_R place5152 (.A(_00112_),
    .Y(net5152));
 BUFx3_ASAP7_75t_R place5153 (.A(_00113_),
    .Y(net5153));
 BUFx3_ASAP7_75t_R place5154 (.A(_00114_),
    .Y(net5154));
 BUFx3_ASAP7_75t_R place5155 (.A(_00115_),
    .Y(net5155));
 BUFx3_ASAP7_75t_R place5156 (.A(_00116_),
    .Y(net5156));
 BUFx3_ASAP7_75t_R place5157 (.A(_00117_),
    .Y(net5157));
 BUFx3_ASAP7_75t_R place5158 (.A(_00118_),
    .Y(net5158));
 BUFx3_ASAP7_75t_R place5162 (.A(_00123_),
    .Y(net5162));
 BUFx3_ASAP7_75t_R place5159 (.A(_00120_),
    .Y(net5159));
 BUFx3_ASAP7_75t_R place5160 (.A(_00121_),
    .Y(net5160));
 BUFx3_ASAP7_75t_R place5161 (.A(_00122_),
    .Y(net5161));
 BUFx3_ASAP7_75t_R place5163 (.A(_00535_),
    .Y(net5163));
 BUFx3_ASAP7_75t_R place5170 (.A(_00133_),
    .Y(net5170));
 BUFx3_ASAP7_75t_R place5164 (.A(_00124_),
    .Y(net5164));
 BUFx3_ASAP7_75t_R place5165 (.A(_00125_),
    .Y(net5165));
 BUFx3_ASAP7_75t_R place5166 (.A(_00127_),
    .Y(net5166));
 BUFx3_ASAP7_75t_R place5167 (.A(_00129_),
    .Y(net5167));
 BUFx3_ASAP7_75t_R place5168 (.A(_00130_),
    .Y(net5168));
 BUFx3_ASAP7_75t_R place5169 (.A(_00131_),
    .Y(net5169));
 BUFx3_ASAP7_75t_R place5171 (.A(_00534_),
    .Y(net5171));
 BUFx3_ASAP7_75t_R place5172 (.A(_00135_),
    .Y(net5172));
 BUFx3_ASAP7_75t_R place5174 (.A(_00138_),
    .Y(net5174));
 BUFx3_ASAP7_75t_R place5175 (.A(_00059_),
    .Y(net5175));
 BUFx3_ASAP7_75t_R place5176 (.A(_00058_),
    .Y(net5176));
 BUFx3_ASAP7_75t_R place5177 (.A(_00139_),
    .Y(net5177));
 BUFx3_ASAP7_75t_R place5178 (.A(_00140_),
    .Y(net5178));
 BUFx3_ASAP7_75t_R place5179 (.A(net5772),
    .Y(net5179));
 BUFx3_ASAP7_75t_R place5180 (.A(_00141_),
    .Y(net5180));
 BUFx3_ASAP7_75t_R place5181 (.A(_00142_),
    .Y(net5181));
 BUFx3_ASAP7_75t_R place5182 (.A(_00143_),
    .Y(net5182));
 BUFx3_ASAP7_75t_R place5183 (.A(_00144_),
    .Y(net5183));
 BUFx3_ASAP7_75t_R place5184 (.A(_00145_),
    .Y(net5184));
 BUFx3_ASAP7_75t_R place5185 (.A(_00146_),
    .Y(net5185));
 BUFx3_ASAP7_75t_R place5186 (.A(_00147_),
    .Y(net5186));
 BUFx3_ASAP7_75t_R place5187 (.A(_00148_),
    .Y(net5187));
 BUFx3_ASAP7_75t_R place5188 (.A(_00149_),
    .Y(net5188));
 BUFx3_ASAP7_75t_R place5189 (.A(_00523_),
    .Y(net5189));
 BUFx3_ASAP7_75t_R place5191 (.A(_00152_),
    .Y(net5191));
 BUFx3_ASAP7_75t_R place5192 (.A(_00153_),
    .Y(net5192));
 BUFx3_ASAP7_75t_R place5193 (.A(_00154_),
    .Y(net5193));
 BUFx3_ASAP7_75t_R place5194 (.A(_00155_),
    .Y(net5194));
 BUFx3_ASAP7_75t_R place5195 (.A(_00159_),
    .Y(net5195));
 BUFx3_ASAP7_75t_R place5196 (.A(_00160_),
    .Y(net5196));
 BUFx3_ASAP7_75t_R place5197 (.A(_00162_),
    .Y(net5197));
 BUFx3_ASAP7_75t_R place5198 (.A(_00336_),
    .Y(net5198));
 BUFx3_ASAP7_75t_R place5199 (.A(_00055_),
    .Y(net5199));
 BUFx3_ASAP7_75t_R place5201 (.A(_00335_),
    .Y(net5201));
 BUFx3_ASAP7_75t_R place5202 (.A(_00334_),
    .Y(net5202));
 BUFx3_ASAP7_75t_R place5203 (.A(_00333_),
    .Y(net5203));
 BUFx3_ASAP7_75t_R place5204 (.A(_00163_),
    .Y(net5204));
 BUFx3_ASAP7_75t_R place5205 (.A(_00331_),
    .Y(net5205));
 BUFx3_ASAP7_75t_R place5211 (.A(_00553_),
    .Y(net5211));
 BUFx3_ASAP7_75t_R place5206 (.A(_00329_),
    .Y(net5206));
 BUFx3_ASAP7_75t_R place5207 (.A(_00164_),
    .Y(net5207));
 BUFx3_ASAP7_75t_R place5208 (.A(_00165_),
    .Y(net5208));
 BUFx3_ASAP7_75t_R place5209 (.A(_00166_),
    .Y(net5209));
 BUFx3_ASAP7_75t_R place5210 (.A(_00169_),
    .Y(net5210));
 BUFx3_ASAP7_75t_R place5212 (.A(_00046_),
    .Y(net5212));
 BUFx3_ASAP7_75t_R place5227 (.A(_00189_),
    .Y(net5227));
 BUFx3_ASAP7_75t_R place5213 (.A(_00327_),
    .Y(net5213));
 BUFx3_ASAP7_75t_R place5214 (.A(_00326_),
    .Y(net5214));
 BUFx3_ASAP7_75t_R place5215 (.A(_00177_),
    .Y(net5215));
 BUFx3_ASAP7_75t_R place5216 (.A(_00178_),
    .Y(net5216));
 BUFx3_ASAP7_75t_R place5217 (.A(_00179_),
    .Y(net5217));
 BUFx3_ASAP7_75t_R place5218 (.A(_00181_),
    .Y(net5218));
 BUFx3_ASAP7_75t_R place5219 (.A(_00182_),
    .Y(net5219));
 BUFx3_ASAP7_75t_R place5220 (.A(_00183_),
    .Y(net5220));
 BUFx3_ASAP7_75t_R place5221 (.A(_00024_),
    .Y(net5221));
 BUFx3_ASAP7_75t_R place5222 (.A(_00184_),
    .Y(net5222));
 BUFx3_ASAP7_75t_R place5223 (.A(_00185_),
    .Y(net5223));
 BUFx3_ASAP7_75t_R place5224 (.A(_00186_),
    .Y(net5224));
 BUFx3_ASAP7_75t_R place5225 (.A(_00187_),
    .Y(net5225));
 BUFx3_ASAP7_75t_R place5226 (.A(_00188_),
    .Y(net5226));
 BUFx3_ASAP7_75t_R place5229 (.A(_00192_),
    .Y(net5229));
 BUFx3_ASAP7_75t_R place5230 (.A(_00193_),
    .Y(net5230));
 BUFx3_ASAP7_75t_R place5231 (.A(_00194_),
    .Y(net5231));
 BUFx3_ASAP7_75t_R place5232 (.A(_00195_),
    .Y(net5232));
 BUFx3_ASAP7_75t_R place5233 (.A(_00196_),
    .Y(net5233));
 BUFx3_ASAP7_75t_R place5234 (.A(_00197_),
    .Y(net5234));
 BUFx3_ASAP7_75t_R place5237 (.A(_00200_),
    .Y(net5237));
 BUFx3_ASAP7_75t_R place5238 (.A(_00201_),
    .Y(net5238));
 BUFx3_ASAP7_75t_R place5239 (.A(_00202_),
    .Y(net5239));
 BUFx3_ASAP7_75t_R place5240 (.A(_00203_),
    .Y(net5240));
 BUFx3_ASAP7_75t_R place5253 (.A(_00224_),
    .Y(net5253));
 BUFx3_ASAP7_75t_R place5241 (.A(_00549_),
    .Y(net5241));
 BUFx3_ASAP7_75t_R place5242 (.A(_00205_),
    .Y(net5242));
 BUFx3_ASAP7_75t_R place5251 (.A(_00061_),
    .Y(net5251));
 BUFx3_ASAP7_75t_R place5243 (.A(_00208_),
    .Y(net5243));
 BUFx3_ASAP7_75t_R place5244 (.A(_00209_),
    .Y(net5244));
 BUFx3_ASAP7_75t_R place5245 (.A(_00210_),
    .Y(net5245));
 BUFx3_ASAP7_75t_R place5246 (.A(_00212_),
    .Y(net5246));
 BUFx3_ASAP7_75t_R place5247 (.A(_00213_),
    .Y(net5247));
 BUFx3_ASAP7_75t_R place5248 (.A(_00214_),
    .Y(net5248));
 BUFx3_ASAP7_75t_R place5249 (.A(_00548_),
    .Y(net5249));
 BUFx3_ASAP7_75t_R place5250 (.A(_00215_),
    .Y(net5250));
 BUFx3_ASAP7_75t_R place5252 (.A(_00062_),
    .Y(net5252));
 BUFx3_ASAP7_75t_R place5255 (.A(_00065_),
    .Y(net5255));
 BUFx3_ASAP7_75t_R place5256 (.A(_00225_),
    .Y(net5256));
 BUFx3_ASAP7_75t_R place5257 (.A(_00226_),
    .Y(net5257));
 BUFx3_ASAP7_75t_R place5258 (.A(_00227_),
    .Y(net5258));
 BUFx3_ASAP7_75t_R place5259 (.A(_00067_),
    .Y(net5259));
 BUFx3_ASAP7_75t_R place5261 (.A(_00057_),
    .Y(net5261));
 BUFx3_ASAP7_75t_R place5262 (.A(_00488_),
    .Y(net5262));
 BUFx3_ASAP7_75t_R place5263 (.A(_00481_),
    .Y(net5263));
 BUFx3_ASAP7_75t_R place5264 (.A(_00480_),
    .Y(net5264));
 BUFx3_ASAP7_75t_R place5265 (.A(_00228_),
    .Y(net5265));
 BUFx3_ASAP7_75t_R place5266 (.A(_00229_),
    .Y(net5266));
 BUFx3_ASAP7_75t_R place5267 (.A(_00230_),
    .Y(net5267));
 BUFx3_ASAP7_75t_R place5268 (.A(_00231_),
    .Y(net5268));
 BUFx3_ASAP7_75t_R place5269 (.A(_00232_),
    .Y(net5269));
 BUFx3_ASAP7_75t_R place5270 (.A(_00233_),
    .Y(net5270));
 BUFx3_ASAP7_75t_R place5271 (.A(_00234_),
    .Y(net5271));
 BUFx3_ASAP7_75t_R place5272 (.A(_00235_),
    .Y(net5272));
 BUFx3_ASAP7_75t_R place5273 (.A(_00396_),
    .Y(net5273));
 BUFx3_ASAP7_75t_R place5274 (.A(_00237_),
    .Y(net5274));
 BUFx3_ASAP7_75t_R place5275 (.A(_00238_),
    .Y(net5275));
 BUFx3_ASAP7_75t_R place5276 (.A(_00239_),
    .Y(net5276));
 BUFx3_ASAP7_75t_R place5277 (.A(_00240_),
    .Y(net5277));
 BUFx3_ASAP7_75t_R place5282 (.A(_00244_),
    .Y(net5282));
 BUFx3_ASAP7_75t_R place5278 (.A(_00241_),
    .Y(net5278));
 BUFx3_ASAP7_75t_R place5279 (.A(_00242_),
    .Y(net5279));
 BUFx3_ASAP7_75t_R place5280 (.A(_00243_),
    .Y(net5280));
 BUFx3_ASAP7_75t_R place5281 (.A(_00365_),
    .Y(net5281));
 BUFx3_ASAP7_75t_R place5284 (.A(_00246_),
    .Y(net5284));
 BUFx3_ASAP7_75t_R place5285 (.A(_00247_),
    .Y(net5285));
 BUFx3_ASAP7_75t_R place5286 (.A(_00248_),
    .Y(net5286));
 BUFx3_ASAP7_75t_R place5288 (.A(_00250_),
    .Y(net5288));
 BUFx3_ASAP7_75t_R place5290 (.A(_00252_),
    .Y(net5290));
 BUFx3_ASAP7_75t_R place5293 (.A(_00255_),
    .Y(net5293));
 BUFx3_ASAP7_75t_R place5294 (.A(_00256_),
    .Y(net5294));
 BUFx3_ASAP7_75t_R place5295 (.A(_00257_),
    .Y(net5295));
 BUFx3_ASAP7_75t_R place5296 (.A(_00259_),
    .Y(net5296));
 BUFx3_ASAP7_75t_R place5297 (.A(_00260_),
    .Y(net5297));
 BUFx3_ASAP7_75t_R place5299 (.A(_00263_),
    .Y(net5299));
 BUFx3_ASAP7_75t_R place5298 (.A(_00262_),
    .Y(net5298));
 BUFx3_ASAP7_75t_R place5301 (.A(_00265_),
    .Y(net5301));
 BUFx3_ASAP7_75t_R place5302 (.A(_00266_),
    .Y(net5302));
 BUFx3_ASAP7_75t_R place5303 (.A(_00267_),
    .Y(net5303));
 BUFx3_ASAP7_75t_R place5304 (.A(_00268_),
    .Y(net5304));
 BUFx3_ASAP7_75t_R place5305 (.A(_00269_),
    .Y(net5305));
 BUFx3_ASAP7_75t_R place5306 (.A(_00270_),
    .Y(net5306));
 BUFx3_ASAP7_75t_R place5307 (.A(_00271_),
    .Y(net5307));
 BUFx3_ASAP7_75t_R place5308 (.A(_00272_),
    .Y(net5308));
 BUFx3_ASAP7_75t_R place5309 (.A(_00273_),
    .Y(net5309));
 BUFx3_ASAP7_75t_R place5310 (.A(_00274_),
    .Y(net5310));
 BUFx3_ASAP7_75t_R place5311 (.A(_00275_),
    .Y(net5311));
 BUFx3_ASAP7_75t_R place5312 (.A(_00276_),
    .Y(net5312));
 BUFx3_ASAP7_75t_R place5313 (.A(_00277_),
    .Y(net5313));
 BUFx3_ASAP7_75t_R place5314 (.A(_00278_),
    .Y(net5314));
 BUFx3_ASAP7_75t_R place5315 (.A(_00279_),
    .Y(net5315));
 BUFx3_ASAP7_75t_R place5316 (.A(_00280_),
    .Y(net5316));
 BUFx3_ASAP7_75t_R place5317 (.A(_00281_),
    .Y(net5317));
 BUFx3_ASAP7_75t_R place5318 (.A(_00282_),
    .Y(net5318));
 BUFx3_ASAP7_75t_R place5319 (.A(_00283_),
    .Y(net5319));
 BUFx3_ASAP7_75t_R place5320 (.A(_00286_),
    .Y(net5320));
 BUFx3_ASAP7_75t_R place5321 (.A(_00287_),
    .Y(net5321));
 BUFx3_ASAP7_75t_R place5322 (.A(_00288_),
    .Y(net5322));
 BUFx3_ASAP7_75t_R place5323 (.A(_00289_),
    .Y(net5323));
 BUFx3_ASAP7_75t_R place5324 (.A(_00290_),
    .Y(net5324));
 BUFx3_ASAP7_75t_R place5325 (.A(_00291_),
    .Y(net5325));
 BUFx3_ASAP7_75t_R place5326 (.A(_00292_),
    .Y(net5326));
 BUFx3_ASAP7_75t_R place5328 (.A(_00294_),
    .Y(net5328));
 BUFx3_ASAP7_75t_R place5329 (.A(_00068_),
    .Y(net5329));
 BUFx3_ASAP7_75t_R place5331 (.A(_00324_),
    .Y(net5331));
 BUFx3_ASAP7_75t_R place5332 (.A(_00323_),
    .Y(net5332));
 BUFx3_ASAP7_75t_R place5360 (.A(_06525_),
    .Y(net5360));
 BUFx3_ASAP7_75t_R place5333 (.A(_00295_),
    .Y(net5333));
 BUFx3_ASAP7_75t_R place5334 (.A(_00296_),
    .Y(net5334));
 BUFx3_ASAP7_75t_R place5335 (.A(_00297_),
    .Y(net5335));
 BUFx3_ASAP7_75t_R place5346 (.A(_00306_),
    .Y(net5346));
 BUFx3_ASAP7_75t_R place5336 (.A(_00476_),
    .Y(net5336));
 BUFx3_ASAP7_75t_R place5337 (.A(_00475_),
    .Y(net5337));
 BUFx3_ASAP7_75t_R place5338 (.A(_00299_),
    .Y(net5338));
 BUFx3_ASAP7_75t_R place5339 (.A(_00300_),
    .Y(net5339));
 BUFx3_ASAP7_75t_R place5340 (.A(_00301_),
    .Y(net5340));
 BUFx3_ASAP7_75t_R place5341 (.A(_00321_),
    .Y(net5341));
 BUFx3_ASAP7_75t_R place5342 (.A(_00320_),
    .Y(net5342));
 BUFx3_ASAP7_75t_R place5343 (.A(_00302_),
    .Y(net5343));
 BUFx3_ASAP7_75t_R place5344 (.A(_00303_),
    .Y(net5344));
 BUFx3_ASAP7_75t_R place5345 (.A(_00304_),
    .Y(net5345));
 BUFx3_ASAP7_75t_R place5347 (.A(_00307_),
    .Y(net5347));
 BUFx6f_ASAP7_75t_R place5359 (.A(net5358),
    .Y(net5359));
 BUFx3_ASAP7_75t_R place5348 (.A(_00308_),
    .Y(net5348));
 BUFx3_ASAP7_75t_R place5349 (.A(_00069_),
    .Y(net5349));
 BUFx3_ASAP7_75t_R place5350 (.A(_00309_),
    .Y(net5350));
 BUFx3_ASAP7_75t_R place5351 (.A(_00310_),
    .Y(net5351));
 BUFx3_ASAP7_75t_R place5352 (.A(_00311_),
    .Y(net5352));
 BUFx3_ASAP7_75t_R place5353 (.A(_00312_),
    .Y(net5353));
 BUFx3_ASAP7_75t_R place5354 (.A(_00313_),
    .Y(net5354));
 BUFx3_ASAP7_75t_R place5355 (.A(_00314_),
    .Y(net5355));
 BUFx3_ASAP7_75t_R place5356 (.A(_00544_),
    .Y(net5356));
 BUFx3_ASAP7_75t_R place5357 (.A(_00543_),
    .Y(net5357));
 BUFx3_ASAP7_75t_R place5358 (.A(_06525_),
    .Y(net5358));
 BUFx24_ASAP7_75t_R clkbuf_leaf_2_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_2_clk));
 BUFx3_ASAP7_75t_R place5363 (.A(net211),
    .Y(net5363));
 BUFx3_ASAP7_75t_R place5362 (.A(net211),
    .Y(net5362));
 BUFx3_ASAP7_75t_R place2753 (.A(_04132_),
    .Y(net2753));
 BUFx3_ASAP7_75t_R place2757 (.A(_04088_),
    .Y(net2757));
 BUFx3_ASAP7_75t_R place2759 (.A(_06414_),
    .Y(net2759));
 BUFx3_ASAP7_75t_R place2761 (.A(_05303_),
    .Y(net2761));
 BUFx3_ASAP7_75t_R place2763 (.A(_04084_),
    .Y(net2763));
 BUFx3_ASAP7_75t_R place2764 (.A(_04084_),
    .Y(net2764));
 BUFx6f_ASAP7_75t_R place2766 (.A(net2765),
    .Y(net2766));
 BUFx3_ASAP7_75t_R place2775 (.A(net2774),
    .Y(net2775));
 BUFx3_ASAP7_75t_R place2780 (.A(_04072_),
    .Y(net2780));
 BUFx3_ASAP7_75t_R place2781 (.A(_06436_),
    .Y(net2781));
 BUFx3_ASAP7_75t_R place2787 (.A(_04102_),
    .Y(net2787));
 BUFx3_ASAP7_75t_R place2791 (.A(net2790),
    .Y(net2791));
 BUFx3_ASAP7_75t_R place2792 (.A(_04063_),
    .Y(net2792));
 BUFx3_ASAP7_75t_R place2801 (.A(_04083_),
    .Y(net2801));
 BUFx3_ASAP7_75t_R place2812 (.A(_05289_),
    .Y(net2812));
 BUFx3_ASAP7_75t_R place2818 (.A(_04057_),
    .Y(net2818));
 BUFx3_ASAP7_75t_R place2826 (.A(_04069_),
    .Y(net2826));
 BUFx3_ASAP7_75t_R place2830 (.A(_02359_),
    .Y(net2830));
 BUFx3_ASAP7_75t_R place2837 (.A(_05282_),
    .Y(net2837));
 BUFx3_ASAP7_75t_R place2839 (.A(net5715),
    .Y(net2839));
 BUFx3_ASAP7_75t_R place2844 (.A(_02368_),
    .Y(net2844));
 BUFx3_ASAP7_75t_R place2845 (.A(_02349_),
    .Y(net2845));
 BUFx3_ASAP7_75t_R place2876 (.A(_02348_),
    .Y(net2876));
 BUFx3_ASAP7_75t_R place2879 (.A(_06380_),
    .Y(net2879));
 BUFx3_ASAP7_75t_R place2881 (.A(_06348_),
    .Y(net2881));
 BUFx3_ASAP7_75t_R place2889 (.A(_02298_),
    .Y(net2889));
 BUFx3_ASAP7_75t_R place2890 (.A(_02287_),
    .Y(net2890));
 BUFx3_ASAP7_75t_R place2891 (.A(_02287_),
    .Y(net2891));
 BUFx3_ASAP7_75t_R place2899 (.A(_06338_),
    .Y(net2899));
 BUFx3_ASAP7_75t_R place2913 (.A(_02306_),
    .Y(net2913));
 BUFx3_ASAP7_75t_R place2922 (.A(_04001_),
    .Y(net2922));
 BUFx3_ASAP7_75t_R place2925 (.A(_02263_),
    .Y(net2925));
 BUFx3_ASAP7_75t_R place2935 (.A(_02256_),
    .Y(net2935));
 BUFx3_ASAP7_75t_R place2943 (.A(net2942),
    .Y(net2943));
 BUFx3_ASAP7_75t_R place2945 (.A(_05194_),
    .Y(net2945));
 BUFx3_ASAP7_75t_R place2947 (.A(_03979_),
    .Y(net2947));
 BUFx3_ASAP7_75t_R place2948 (.A(_03971_),
    .Y(net2948));
 BUFx3_ASAP7_75t_R place2958 (.A(_06297_),
    .Y(net2958));
 BUFx3_ASAP7_75t_R place2963 (.A(net2962),
    .Y(net2963));
 BUFx3_ASAP7_75t_R place2967 (.A(_03970_),
    .Y(net2967));
 BUFx3_ASAP7_75t_R place3013 (.A(_05148_),
    .Y(net3013));
 BUFx3_ASAP7_75t_R place3014 (.A(_03951_),
    .Y(net3014));
 BUFx3_ASAP7_75t_R place3059 (.A(_06238_),
    .Y(net3059));
 BUFx3_ASAP7_75t_R place3063 (.A(_03932_),
    .Y(net3063));
 BUFx6f_ASAP7_75t_R place3064 (.A(_03915_),
    .Y(net3064));
 BUFx3_ASAP7_75t_R place3065 (.A(net3064),
    .Y(net3065));
 BUFx3_ASAP7_75t_R place3095 (.A(_05085_),
    .Y(net3095));
 BUFx3_ASAP7_75t_R place3101 (.A(_05118_),
    .Y(net3101));
 BUFx3_ASAP7_75t_R place3118 (.A(_02151_),
    .Y(net3118));
 BUFx3_ASAP7_75t_R place3126 (.A(_03825_),
    .Y(net3126));
 BUFx3_ASAP7_75t_R place3130 (.A(_02125_),
    .Y(net3130));
 BUFx3_ASAP7_75t_R place3131 (.A(net3130),
    .Y(net3131));
 BUFx3_ASAP7_75t_R place3160 (.A(_06180_),
    .Y(net3160));
 BUFx3_ASAP7_75t_R place3161 (.A(_06168_),
    .Y(net3161));
 BUFx3_ASAP7_75t_R place3167 (.A(_03798_),
    .Y(net3167));
 BUFx3_ASAP7_75t_R place3177 (.A(_06129_),
    .Y(net3177));
 BUFx3_ASAP7_75t_R place3195 (.A(_06121_),
    .Y(net3195));
 BUFx3_ASAP7_75t_R place3196 (.A(_06121_),
    .Y(net3196));
 BUFx3_ASAP7_75t_R place3197 (.A(net3196),
    .Y(net3197));
 BUFx3_ASAP7_75t_R place3212 (.A(_06133_),
    .Y(net3212));
 BUFx3_ASAP7_75t_R place3229 (.A(_05015_),
    .Y(net3229));
 BUFx3_ASAP7_75t_R place3231 (.A(_03820_),
    .Y(net3231));
 BUFx3_ASAP7_75t_R place3238 (.A(_06126_),
    .Y(net3238));
 BUFx3_ASAP7_75t_R place3242 (.A(_03791_),
    .Y(net3242));
 BUFx3_ASAP7_75t_R place3244 (.A(_02082_),
    .Y(net3244));
 BUFx6f_ASAP7_75t_R place3246 (.A(_02075_),
    .Y(net3246));
 BUFx3_ASAP7_75t_R place3247 (.A(net3246),
    .Y(net3247));
 BUFx3_ASAP7_75t_R place3258 (.A(net3257),
    .Y(net3258));
 BUFx3_ASAP7_75t_R place3265 (.A(_03737_),
    .Y(net3265));
 BUFx3_ASAP7_75t_R place3267 (.A(_02037_),
    .Y(net3267));
 BUFx3_ASAP7_75t_R place3276 (.A(_03736_),
    .Y(net3276));
 BUFx3_ASAP7_75t_R place3325 (.A(_04969_),
    .Y(net3325));
 BUFx3_ASAP7_75t_R place3331 (.A(_03753_),
    .Y(net3331));
 BUFx3_ASAP7_75t_R place3333 (.A(net5678),
    .Y(net3333));
 BUFx3_ASAP7_75t_R place3335 (.A(net3334),
    .Y(net3335));
 BUFx3_ASAP7_75t_R place3459 (.A(_03647_),
    .Y(net3459));
 BUFx3_ASAP7_75t_R place3535 (.A(net5679),
    .Y(net3535));
 BUFx3_ASAP7_75t_R place3548 (.A(_03594_),
    .Y(net3548));
 BUFx3_ASAP7_75t_R place3572 (.A(_04793_),
    .Y(net3572));
 BUFx3_ASAP7_75t_R place3576 (.A(_03585_),
    .Y(net3576));
 BUFx3_ASAP7_75t_R place3590 (.A(_04792_),
    .Y(net3590));
 BUFx3_ASAP7_75t_R place3593 (.A(_03554_),
    .Y(net3593));
 BUFx3_ASAP7_75t_R place3618 (.A(_01807_),
    .Y(net3618));
 BUFx3_ASAP7_75t_R place3623 (.A(_05866_),
    .Y(net3623));
 BUFx3_ASAP7_75t_R place3633 (.A(net3632),
    .Y(net3633));
 BUFx3_ASAP7_75t_R place3635 (.A(_03544_),
    .Y(net3635));
 BUFx3_ASAP7_75t_R place3636 (.A(net3635),
    .Y(net3636));
 BUFx6f_ASAP7_75t_R place3641 (.A(_01811_),
    .Y(net3641));
 BUFx3_ASAP7_75t_R place3646 (.A(net3645),
    .Y(net3646));
 BUFx3_ASAP7_75t_R place3659 (.A(net3658),
    .Y(net3659));
 BUFx3_ASAP7_75t_R place3677 (.A(_01751_),
    .Y(net3677));
 BUFx3_ASAP7_75t_R place3705 (.A(_01754_),
    .Y(net3705));
 BUFx3_ASAP7_75t_R place3707 (.A(_05828_),
    .Y(net3707));
 BUFx3_ASAP7_75t_R place3711 (.A(_03500_),
    .Y(net3711));
 BUFx3_ASAP7_75t_R place3713 (.A(_03471_),
    .Y(net3713));
 BUFx3_ASAP7_75t_R place3714 (.A(_01753_),
    .Y(net3714));
 BUFx3_ASAP7_75t_R place3715 (.A(net5764),
    .Y(net3715));
 BUFx3_ASAP7_75t_R place3725 (.A(_01745_),
    .Y(net3725));
 BUFx3_ASAP7_75t_R place3727 (.A(_01743_),
    .Y(net3727));
 BUFx6f_ASAP7_75t_R place3734 (.A(_05798_),
    .Y(net3734));
 BUFx3_ASAP7_75t_R place3754 (.A(net5757),
    .Y(net3754));
 BUFx3_ASAP7_75t_R place3755 (.A(_01716_),
    .Y(net3755));
 BUFx3_ASAP7_75t_R place3770 (.A(_03433_),
    .Y(net3770));
 BUFx3_ASAP7_75t_R place3776 (.A(_01683_),
    .Y(net3776));
 BUFx3_ASAP7_75t_R place3788 (.A(net5975),
    .Y(net3788));
 BUFx3_ASAP7_75t_R place3790 (.A(_03431_),
    .Y(net3790));
 BUFx3_ASAP7_75t_R place3793 (.A(_01703_),
    .Y(net3793));
 BUFx3_ASAP7_75t_R place3808 (.A(_05753_),
    .Y(net3808));
 BUFx3_ASAP7_75t_R place3810 (.A(_04667_),
    .Y(net3810));
 BUFx3_ASAP7_75t_R place3812 (.A(net3811),
    .Y(net3812));
 BUFx3_ASAP7_75t_R place3821 (.A(_05714_),
    .Y(net3821));
 BUFx3_ASAP7_75t_R place3822 (.A(net5613),
    .Y(net3822));
 BUFx3_ASAP7_75t_R place3826 (.A(net3825),
    .Y(net3826));
 BUFx3_ASAP7_75t_R place3922 (.A(_01626_),
    .Y(net3922));
 BUFx3_ASAP7_75t_R place3927 (.A(_01566_),
    .Y(net3927));
 BUFx6f_ASAP7_75t_R place3931 (.A(net3930),
    .Y(net3931));
 BUFx3_ASAP7_75t_R place3934 (.A(_01615_),
    .Y(net3934));
 BUFx3_ASAP7_75t_R place3940 (.A(_04581_),
    .Y(net3940));
 BUFx3_ASAP7_75t_R place3953 (.A(_01585_),
    .Y(net3953));
 BUFx3_ASAP7_75t_R place3983 (.A(_03312_),
    .Y(net3983));
 BUFx3_ASAP7_75t_R place3984 (.A(_03312_),
    .Y(net3984));
 BUFx3_ASAP7_75t_R place3988 (.A(_04504_),
    .Y(net3988));
 BUFx3_ASAP7_75t_R place4041 (.A(net4040),
    .Y(net4041));
 BUFx3_ASAP7_75t_R place4052 (.A(net4051),
    .Y(net4052));
 BUFx3_ASAP7_75t_R place4065 (.A(_05604_),
    .Y(net4065));
 BUFx3_ASAP7_75t_R place4069 (.A(_04677_),
    .Y(net4069));
 BUFx3_ASAP7_75t_R place4075 (.A(net4074),
    .Y(net4075));
 BUFx3_ASAP7_75t_R place4086 (.A(net4085),
    .Y(net4086));
 BUFx3_ASAP7_75t_R place4106 (.A(_06007_),
    .Y(net4106));
 BUFx3_ASAP7_75t_R place4107 (.A(_05917_),
    .Y(net4107));
 BUFx3_ASAP7_75t_R place4125 (.A(_04790_),
    .Y(net4125));
 BUFx3_ASAP7_75t_R place4128 (.A(_04726_),
    .Y(net4128));
 BUFx3_ASAP7_75t_R place4133 (.A(net4132),
    .Y(net4133));
 BUFx3_ASAP7_75t_R place4147 (.A(net4146),
    .Y(net4147));
 BUFx3_ASAP7_75t_R place4157 (.A(net4156),
    .Y(net4157));
 BUFx3_ASAP7_75t_R place4160 (.A(net4159),
    .Y(net4160));
 BUFx6f_ASAP7_75t_R place4162 (.A(_02064_),
    .Y(net4162));
 BUFx3_ASAP7_75t_R place4163 (.A(net4162),
    .Y(net4163));
 BUFx3_ASAP7_75t_R place4167 (.A(net4166),
    .Y(net4167));
 BUFx6f_ASAP7_75t_R place4169 (.A(net4168),
    .Y(net4169));
 BUFx3_ASAP7_75t_R place4181 (.A(net4180),
    .Y(net4181));
 BUFx3_ASAP7_75t_R place4258 (.A(net4257),
    .Y(net4258));
 BUFx3_ASAP7_75t_R place4259 (.A(_05173_),
    .Y(net4259));
 BUFx6f_ASAP7_75t_R place4260 (.A(net4259),
    .Y(net4260));
 BUFx3_ASAP7_75t_R place4261 (.A(net4260),
    .Y(net4261));
 BUFx3_ASAP7_75t_R place4288 (.A(net4286),
    .Y(net4288));
 BUFx3_ASAP7_75t_R place4289 (.A(net4286),
    .Y(net4289));
 BUFx3_ASAP7_75t_R place4290 (.A(net4289),
    .Y(net4290));
 BUFx3_ASAP7_75t_R place4310 (.A(_05477_),
    .Y(net4310));
 BUFx3_ASAP7_75t_R place4342 (.A(net4340),
    .Y(net4342));
 BUFx3_ASAP7_75t_R place4349 (.A(net5607),
    .Y(net4349));
 BUFx3_ASAP7_75t_R place4353 (.A(_04457_),
    .Y(net4353));
 BUFx3_ASAP7_75t_R place4355 (.A(net4354),
    .Y(net4355));
 BUFx3_ASAP7_75t_R place4363 (.A(net4361),
    .Y(net4363));
 BUFx3_ASAP7_75t_R place4397 (.A(net4396),
    .Y(net4397));
 BUFx3_ASAP7_75t_R place4401 (.A(_05472_),
    .Y(net4401));
 BUFx3_ASAP7_75t_R place4402 (.A(_05472_),
    .Y(net4402));
 BUFx3_ASAP7_75t_R place4425 (.A(_03239_),
    .Y(net4425));
 BUFx3_ASAP7_75t_R place4427 (.A(_03217_),
    .Y(net4427));
 BUFx3_ASAP7_75t_R place4430 (.A(_02622_),
    .Y(net4430));
 BUFx3_ASAP7_75t_R place4431 (.A(_02591_),
    .Y(net4431));
 BUFx3_ASAP7_75t_R place4593 (.A(_01186_),
    .Y(net4593));
 BUFx3_ASAP7_75t_R place4594 (.A(_01168_),
    .Y(net4594));
 BUFx3_ASAP7_75t_R place4595 (.A(_01161_),
    .Y(net4595));
 BUFx3_ASAP7_75t_R place4656 (.A(net4655),
    .Y(net4656));
 BUFx6f_ASAP7_75t_R place5049 (.A(_00929_),
    .Y(net5049));
 BUFx3_ASAP7_75t_R place5050 (.A(net5049),
    .Y(net5050));
 BUFx6f_ASAP7_75t_R place5051 (.A(net5049),
    .Y(net5051));
 BUFx6f_ASAP7_75t_R place5052 (.A(net5049),
    .Y(net5052));
 BUFx6f_ASAP7_75t_R place5053 (.A(net5049),
    .Y(net5053));
 BUFx3_ASAP7_75t_R place5054 (.A(net5049),
    .Y(net5054));
 BUFx6f_ASAP7_75t_R place5055 (.A(net5049),
    .Y(net5055));
 BUFx3_ASAP7_75t_R place5059 (.A(_00909_),
    .Y(net5059));
 BUFx3_ASAP7_75t_R place5060 (.A(_00908_),
    .Y(net5060));
 BUFx3_ASAP7_75t_R place5062 (.A(_00903_),
    .Y(net5062));
 BUFx3_ASAP7_75t_R place5063 (.A(_00896_),
    .Y(net5063));
 BUFx3_ASAP7_75t_R place5069 (.A(\u_fft.sched[42] ),
    .Y(net5069));
 BUFx3_ASAP7_75t_R place5088 (.A(_00025_),
    .Y(net5088));
 BUFx3_ASAP7_75t_R place5200 (.A(net5199),
    .Y(net5200));
 BUFx3_ASAP7_75t_R place5228 (.A(_00191_),
    .Y(net5228));
 BUFx3_ASAP7_75t_R place5235 (.A(_00198_),
    .Y(net5235));
 BUFx3_ASAP7_75t_R place5236 (.A(_00199_),
    .Y(net5236));
 BUFx3_ASAP7_75t_R place5254 (.A(_00063_),
    .Y(net5254));
 BUFx3_ASAP7_75t_R place5260 (.A(net5259),
    .Y(net5260));
 BUFx3_ASAP7_75t_R place5283 (.A(_00245_),
    .Y(net5283));
 BUFx3_ASAP7_75t_R place5287 (.A(_00249_),
    .Y(net5287));
 BUFx3_ASAP7_75t_R place5289 (.A(_00251_),
    .Y(net5289));
 BUFx3_ASAP7_75t_R place5291 (.A(_00253_),
    .Y(net5291));
 BUFx3_ASAP7_75t_R place5292 (.A(_00254_),
    .Y(net5292));
 BUFx3_ASAP7_75t_R place5300 (.A(_00264_),
    .Y(net5300));
 BUFx3_ASAP7_75t_R place5327 (.A(_00293_),
    .Y(net5327));
 BUFx3_ASAP7_75t_R place5330 (.A(net5329),
    .Y(net5330));
 BUFx6f_ASAP7_75t_R place5361 (.A(net5360),
    .Y(net5361));
 BUFx24_ASAP7_75t_R clkbuf_leaf_3_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_3_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_4_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_4_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_5_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_5_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_6_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_6_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_7_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_7_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_8_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_8_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_9_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_9_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_10_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_10_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_11_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_11_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_12_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_12_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_13_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_13_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_14_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_14_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_15_clk (.A(clknet_1_1__leaf_clk),
    .Y(clknet_leaf_15_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_16_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_16_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_17_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_17_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_18_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_18_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_19_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_19_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_20_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_20_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_21_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_21_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_22_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_22_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_23_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_23_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_24_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_24_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_25_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_25_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_26_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_26_clk));
 BUFx24_ASAP7_75t_R clkbuf_leaf_27_clk (.A(clknet_1_0__leaf_clk),
    .Y(clknet_leaf_27_clk));
 BUFx24_ASAP7_75t_R clkbuf_0_clk (.A(clk),
    .Y(clknet_0_clk));
 BUFx24_ASAP7_75t_R clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Y(clknet_1_0__leaf_clk));
 BUFx24_ASAP7_75t_R clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Y(clknet_1_1__leaf_clk));
 BUFx12_ASAP7_75t_R clkload0 (.A(clknet_leaf_0_clk));
 INVx3_ASAP7_75t_R clkload1 (.A(clknet_leaf_16_clk));
 BUFx12_ASAP7_75t_R clkload2 (.A(clknet_leaf_17_clk));
 BUFx12_ASAP7_75t_R clkload3 (.A(clknet_leaf_18_clk));
 INVx3_ASAP7_75t_R clkload4 (.A(clknet_leaf_19_clk));
 BUFx2_ASAP7_75t_R clkload5 (.A(clknet_leaf_20_clk));
 BUFx2_ASAP7_75t_R clkload6 (.A(clknet_leaf_21_clk));
 BUFx4f_ASAP7_75t_R clkload7 (.A(clknet_leaf_22_clk));
 BUFx2_ASAP7_75t_R clkload8 (.A(clknet_leaf_23_clk));
 BUFx4f_ASAP7_75t_R clkload9 (.A(clknet_leaf_24_clk));
 INVx3_ASAP7_75t_R clkload10 (.A(clknet_leaf_25_clk));
 INVx3_ASAP7_75t_R clkload11 (.A(clknet_leaf_26_clk));
 INVx6_ASAP7_75t_R clkload12 (.A(clknet_leaf_27_clk));
 INVx5_ASAP7_75t_R clkload13 (.A(clknet_leaf_1_clk));
 BUFx12_ASAP7_75t_R clkload14 (.A(clknet_leaf_4_clk));
 BUFx4f_ASAP7_75t_R clkload15 (.A(clknet_leaf_5_clk));
 BUFx12_ASAP7_75t_R clkload16 (.A(clknet_leaf_6_clk));
 BUFx4f_ASAP7_75t_R clkload17 (.A(clknet_leaf_7_clk));
 BUFx24_ASAP7_75t_R clkload18 (.A(clknet_leaf_8_clk));
 INVx8_ASAP7_75t_R clkload19 (.A(clknet_leaf_9_clk));
 INVx5_ASAP7_75t_R clkload20 (.A(clknet_leaf_10_clk));
 BUFx24_ASAP7_75t_R clkload21 (.A(clknet_leaf_11_clk));
 INVx3_ASAP7_75t_R clkload22 (.A(clknet_leaf_12_clk));
 INVx8_ASAP7_75t_R clkload23 (.A(clknet_leaf_13_clk));
 BUFx2_ASAP7_75t_R clkload24 (.A(clknet_leaf_14_clk));
 CKINVDCx10_ASAP7_75t_R clkload25 (.A(clknet_leaf_15_clk));
 BUFx3_ASAP7_75t_R rebuffer5364 (.A(_00458_),
    .Y(net5364));
 BUFx3_ASAP7_75t_R rebuffer5365 (.A(net5364),
    .Y(net5365));
 BUFx3_ASAP7_75t_R rebuffer5366 (.A(_00418_),
    .Y(net5366));
 BUFx3_ASAP7_75t_R rebuffer5367 (.A(_00438_),
    .Y(net5367));
 BUFx3_ASAP7_75t_R rebuffer5368 (.A(_01284_),
    .Y(net5368));
 BUFx3_ASAP7_75t_R rebuffer5369 (.A(_00416_),
    .Y(net5369));
 BUFx3_ASAP7_75t_R rebuffer5370 (.A(_01318_),
    .Y(net5370));
 BUFx3_ASAP7_75t_R rebuffer5371 (.A(_01058_),
    .Y(net5371));
 BUFx6f_ASAP7_75t_R rebuffer5372 (.A(net5419),
    .Y(net5372));
 BUFx6f_ASAP7_75t_R rebuffer5373 (.A(_02229_),
    .Y(net5373));
 BUFx3_ASAP7_75t_R rebuffer5374 (.A(net5373),
    .Y(net5374));
 BUFx3_ASAP7_75t_R rebuffer5375 (.A(_00408_),
    .Y(net5375));
 BUFx3_ASAP7_75t_R rebuffer5376 (.A(net5375),
    .Y(net5376));
 BUFx6f_ASAP7_75t_R rebuffer5377 (.A(_01051_),
    .Y(net5377));
 BUFx3_ASAP7_75t_R rebuffer5378 (.A(_00439_),
    .Y(net5378));
 BUFx3_ASAP7_75t_R rebuffer5379 (.A(_01340_),
    .Y(net5379));
 BUFx3_ASAP7_75t_R rebuffer5380 (.A(_01357_),
    .Y(net5380));
 BUFx6f_ASAP7_75t_R rebuffer5381 (.A(_01159_),
    .Y(net5381));
 BUFx3_ASAP7_75t_R rebuffer5382 (.A(_02164_),
    .Y(net5382));
 BUFx3_ASAP7_75t_R rebuffer5383 (.A(_01809_),
    .Y(net5383));
 BUFx3_ASAP7_75t_R rebuffer5384 (.A(_01279_),
    .Y(net5384));
 BUFx6f_ASAP7_75t_R rebuffer5385 (.A(_01422_),
    .Y(net5385));
 BUFx3_ASAP7_75t_R rebuffer5386 (.A(_01501_),
    .Y(net5386));
 BUFx3_ASAP7_75t_R rebuffer5387 (.A(_02039_),
    .Y(net5387));
 BUFx3_ASAP7_75t_R rebuffer5388 (.A(_01909_),
    .Y(net5388));
 BUFx3_ASAP7_75t_R rebuffer5389 (.A(_01899_),
    .Y(net5389));
 BUFx3_ASAP7_75t_R rebuffer5390 (.A(_01899_),
    .Y(net5390));
 BUFx3_ASAP7_75t_R rebuffer5391 (.A(_02293_),
    .Y(net5391));
 BUFx3_ASAP7_75t_R rebuffer5392 (.A(_02071_),
    .Y(net5392));
 BUFx3_ASAP7_75t_R rebuffer5393 (.A(net4767),
    .Y(net5393));
 BUFx6f_ASAP7_75t_R clone5394 (.A(_02387_),
    .Y(net5394));
 BUFx3_ASAP7_75t_R rebuffer5395 (.A(_00076_),
    .Y(net5395));
 BUFx3_ASAP7_75t_R rebuffer5396 (.A(_02130_),
    .Y(net5396));
 BUFx6f_ASAP7_75t_R rebuffer5397 (.A(_02163_),
    .Y(net5397));
 BUFx3_ASAP7_75t_R rebuffer5398 (.A(_02300_),
    .Y(net5398));
 BUFx3_ASAP7_75t_R rebuffer5399 (.A(_01673_),
    .Y(net5399));
 BUFx3_ASAP7_75t_R rebuffer5400 (.A(net5399),
    .Y(net5400));
 BUFx6f_ASAP7_75t_R rebuffer5401 (.A(_01829_),
    .Y(net5401));
 BUFx3_ASAP7_75t_R rebuffer5402 (.A(_01231_),
    .Y(net5402));
 BUFx6f_ASAP7_75t_R rebuffer5403 (.A(_01311_),
    .Y(net5403));
 BUFx3_ASAP7_75t_R rebuffer5404 (.A(_01311_),
    .Y(net5404));
 BUFx12f_ASAP7_75t_R clone5418 (.A(net5903),
    .Y(net5418));
 BUFx6f_ASAP7_75t_R rebuffer5419 (.A(_02523_),
    .Y(net5419));
 BUFx3_ASAP7_75t_R rebuffer5420 (.A(_02384_),
    .Y(net5420));
 BUFx6f_ASAP7_75t_R rebuffer5421 (.A(_02255_),
    .Y(net5421));
 BUFx3_ASAP7_75t_R rebuffer5422 (.A(_02013_),
    .Y(net5422));
 BUFx3_ASAP7_75t_R rebuffer5423 (.A(_01941_),
    .Y(net5423));
 BUFx6f_ASAP7_75t_R rebuffer5424 (.A(_01932_),
    .Y(net5424));
 BUFx3_ASAP7_75t_R rebuffer5425 (.A(_01444_),
    .Y(net5425));
 BUFx3_ASAP7_75t_R rebuffer5426 (.A(_01449_),
    .Y(net5426));
 BUFx3_ASAP7_75t_R rebuffer5427 (.A(_01323_),
    .Y(net5427));
 BUFx3_ASAP7_75t_R rebuffer5428 (.A(_01417_),
    .Y(net5428));
 BUFx3_ASAP7_75t_R rebuffer5429 (.A(_01259_),
    .Y(net5429));
 BUFx3_ASAP7_75t_R rebuffer5430 (.A(_01594_),
    .Y(net5430));
 BUFx3_ASAP7_75t_R rebuffer5431 (.A(net5902),
    .Y(net5431));
 BUFx6f_ASAP7_75t_R rebuffer5432 (.A(_01052_),
    .Y(net5432));
 BUFx3_ASAP7_75t_R rebuffer5433 (.A(_01308_),
    .Y(net5433));
 BUFx3_ASAP7_75t_R rebuffer5434 (.A(\u_window_buffer.read_ptr[14] ),
    .Y(net5434));
 BUFx3_ASAP7_75t_R rebuffer5435 (.A(net4765),
    .Y(net5435));
 BUFx3_ASAP7_75t_R rebuffer5436 (.A(net4771),
    .Y(net5436));
 BUFx3_ASAP7_75t_R rebuffer5437 (.A(_01667_),
    .Y(net5437));
 BUFx3_ASAP7_75t_R rebuffer5438 (.A(_01713_),
    .Y(net5438));
 BUFx6f_ASAP7_75t_R rebuffer5439 (.A(_02014_),
    .Y(net5439));
 BUFx3_ASAP7_75t_R rebuffer5440 (.A(_02083_),
    .Y(net5440));
 BUFx3_ASAP7_75t_R rebuffer5441 (.A(_02083_),
    .Y(net5441));
 BUFx3_ASAP7_75t_R rebuffer5442 (.A(_02031_),
    .Y(net5442));
 BUFx3_ASAP7_75t_R rebuffer5443 (.A(_02061_),
    .Y(net5443));
 BUFx3_ASAP7_75t_R rebuffer5444 (.A(_01999_),
    .Y(net5444));
 BUFx3_ASAP7_75t_R rebuffer5445 (.A(_02275_),
    .Y(net5445));
 BUFx3_ASAP7_75t_R rebuffer5446 (.A(_02275_),
    .Y(net5446));
 BUFx3_ASAP7_75t_R rebuffer5447 (.A(_02279_),
    .Y(net5447));
 BUFx3_ASAP7_75t_R rebuffer5448 (.A(_02277_),
    .Y(net5448));
 BUFx3_ASAP7_75t_R rebuffer5449 (.A(_02165_),
    .Y(net5449));
 BUFx3_ASAP7_75t_R rebuffer5450 (.A(_01955_),
    .Y(net5450));
 BUFx3_ASAP7_75t_R rebuffer5451 (.A(net5887),
    .Y(net5451));
 BUFx3_ASAP7_75t_R rebuffer5452 (.A(_02246_),
    .Y(net5452));
 BUFx3_ASAP7_75t_R rebuffer5453 (.A(_02246_),
    .Y(net5453));
 BUFx3_ASAP7_75t_R rebuffer5454 (.A(_02070_),
    .Y(net5454));
 BUFx3_ASAP7_75t_R rebuffer5455 (.A(_01679_),
    .Y(net5455));
 BUFx3_ASAP7_75t_R rebuffer5456 (.A(net3541),
    .Y(net5456));
 BUFx3_ASAP7_75t_R rebuffer5457 (.A(\u_window_buffer.read_ptr[6] ),
    .Y(net5457));
 BUFx3_ASAP7_75t_R rebuffer5458 (.A(_02204_),
    .Y(net5458));
 BUFx6f_ASAP7_75t_R rebuffer5504 (.A(_04329_),
    .Y(net5504));
 BUFx3_ASAP7_75t_R rebuffer5505 (.A(_02342_),
    .Y(net5505));
 BUFx6f_ASAP7_75t_R rebuffer5506 (.A(net2709),
    .Y(net5506));
 BUFx3_ASAP7_75t_R clone5536 (.A(_02524_),
    .Y(net5536));
 BUFx3_ASAP7_75t_R rebuffer5537 (.A(_02318_),
    .Y(net5537));
 BUFx6f_ASAP7_75t_R rebuffer5538 (.A(net5541),
    .Y(net5538));
 BUFx3_ASAP7_75t_R rebuffer5539 (.A(net5541),
    .Y(net5539));
 BUFx6f_ASAP7_75t_R rebuffer5540 (.A(net5541),
    .Y(net5540));
 BUFx6f_ASAP7_75t_R clone5541 (.A(net5590),
    .Y(net5541));
 BUFx3_ASAP7_75t_R rebuffer5585 (.A(_00100_),
    .Y(net5585));
 BUFx3_ASAP7_75t_R rebuffer5590 (.A(net2709),
    .Y(net5590));
 BUFx6f_ASAP7_75t_R clone5591 (.A(_05355_),
    .Y(net5591));
 BUFx6f_ASAP7_75t_R rebuffer5592 (.A(net2709),
    .Y(net5592));
 BUFx6f_ASAP7_75t_R rebuffer5593 (.A(_05776_),
    .Y(net5593));
 BUFx3_ASAP7_75t_R rebuffer5594 (.A(_05776_),
    .Y(net5594));
 BUFx3_ASAP7_75t_R rebuffer5595 (.A(_05890_),
    .Y(net5595));
 BUFx3_ASAP7_75t_R rebuffer5596 (.A(_06038_),
    .Y(net5596));
 BUFx3_ASAP7_75t_R rebuffer5597 (.A(_06260_),
    .Y(net5597));
 BUFx3_ASAP7_75t_R rebuffer5598 (.A(_06397_),
    .Y(net5598));
 BUFx3_ASAP7_75t_R rebuffer5599 (.A(_05836_),
    .Y(net5599));
 BUFx3_ASAP7_75t_R rebuffer5600 (.A(net5601),
    .Y(net5600));
 BUFx3_ASAP7_75t_R rebuffer5601 (.A(_06051_),
    .Y(net5601));
 BUFx3_ASAP7_75t_R rebuffer5602 (.A(_06258_),
    .Y(net5602));
 BUFx3_ASAP7_75t_R rebuffer5603 (.A(_00541_),
    .Y(net5603));
 BUFx3_ASAP7_75t_R rebuffer5604 (.A(_05425_),
    .Y(net5604));
 BUFx3_ASAP7_75t_R rebuffer5605 (.A(_06152_),
    .Y(net5605));
 BUFx3_ASAP7_75t_R rebuffer5606 (.A(_06323_),
    .Y(net5606));
 BUFx3_ASAP7_75t_R rebuffer5607 (.A(_05502_),
    .Y(net5607));
 BUFx3_ASAP7_75t_R rebuffer5608 (.A(_05707_),
    .Y(net5608));
 BUFx3_ASAP7_75t_R rebuffer5609 (.A(_05739_),
    .Y(net5609));
 BUFx3_ASAP7_75t_R rebuffer5610 (.A(_05933_),
    .Y(net5610));
 BUFx3_ASAP7_75t_R rebuffer5611 (.A(_05855_),
    .Y(net5611));
 BUFx3_ASAP7_75t_R rebuffer5612 (.A(_05650_),
    .Y(net5612));
 BUFx3_ASAP7_75t_R rebuffer5613 (.A(_05714_),
    .Y(net5613));
 BUFx3_ASAP7_75t_R rebuffer5614 (.A(_06370_),
    .Y(net5614));
 BUFx3_ASAP7_75t_R rebuffer5615 (.A(_06269_),
    .Y(net5615));
 BUFx3_ASAP7_75t_R rebuffer5616 (.A(_05764_),
    .Y(net5616));
 BUFx3_ASAP7_75t_R rebuffer5617 (.A(net5616),
    .Y(net5617));
 BUFx3_ASAP7_75t_R rebuffer5618 (.A(net5958),
    .Y(net5618));
 BUFx3_ASAP7_75t_R rebuffer5619 (.A(_06100_),
    .Y(net5619));
 BUFx3_ASAP7_75t_R rebuffer5620 (.A(_06332_),
    .Y(net5620));
 BUFx6f_ASAP7_75t_R rebuffer5621 (.A(_06232_),
    .Y(net5621));
 BUFx3_ASAP7_75t_R rebuffer5622 (.A(_06420_),
    .Y(net5622));
 BUFx3_ASAP7_75t_R rebuffer5623 (.A(\u_window_buffer.write_ptr[1] ),
    .Y(net5623));
 BUFx6f_ASAP7_75t_R rebuffer5624 (.A(_06054_),
    .Y(net5624));
 BUFx3_ASAP7_75t_R rebuffer5625 (.A(_06084_),
    .Y(net5625));
 BUFx3_ASAP7_75t_R rebuffer5626 (.A(_06258_),
    .Y(net5626));
 BUFx3_ASAP7_75t_R rebuffer5627 (.A(_06190_),
    .Y(net5627));
 BUFx3_ASAP7_75t_R rebuffer5628 (.A(_06029_),
    .Y(net5628));
 BUFx3_ASAP7_75t_R rebuffer5629 (.A(_05975_),
    .Y(net5629));
 BUFx3_ASAP7_75t_R rebuffer5630 (.A(_06061_),
    .Y(net5630));
 BUFx3_ASAP7_75t_R rebuffer5631 (.A(_06059_),
    .Y(net5631));
 BUFx3_ASAP7_75t_R rebuffer5632 (.A(_06036_),
    .Y(net5632));
 BUFx3_ASAP7_75t_R rebuffer5633 (.A(_06111_),
    .Y(net5633));
 BUFx6f_ASAP7_75t_R rebuffer5634 (.A(_06155_),
    .Y(net5634));
 BUFx3_ASAP7_75t_R rebuffer5635 (.A(net5115),
    .Y(net5635));
 BUFx3_ASAP7_75t_R rebuffer5636 (.A(_06327_),
    .Y(net5636));
 BUFx3_ASAP7_75t_R rebuffer5637 (.A(_06328_),
    .Y(net5637));
 BUFx3_ASAP7_75t_R rebuffer5638 (.A(_05996_),
    .Y(net5638));
 BUFx3_ASAP7_75t_R rebuffer5653 (.A(_06443_),
    .Y(net5653));
 BUFx3_ASAP7_75t_R rebuffer5654 (.A(net3976),
    .Y(net5654));
 BUFx3_ASAP7_75t_R rebuffer5655 (.A(_05620_),
    .Y(net5655));
 BUFx3_ASAP7_75t_R rebuffer5661 (.A(_06469_),
    .Y(net5661));
 BUFx3_ASAP7_75t_R rebuffer5662 (.A(_06466_),
    .Y(net5662));
 BUFx3_ASAP7_75t_R rebuffer5663 (.A(_06196_),
    .Y(net5663));
 BUFx3_ASAP7_75t_R rebuffer5664 (.A(net2825),
    .Y(net5664));
 BUFx3_ASAP7_75t_R rebuffer5665 (.A(_05498_),
    .Y(net5665));
 BUFx3_ASAP7_75t_R rebuffer5666 (.A(net5695),
    .Y(net5666));
 BUFx6f_ASAP7_75t_R rebuffer5667 (.A(_03576_),
    .Y(net5667));
 BUFx3_ASAP7_75t_R rebuffer5668 (.A(_03576_),
    .Y(net5668));
 BUFx3_ASAP7_75t_R rebuffer5669 (.A(net5981),
    .Y(net5669));
 BUFx3_ASAP7_75t_R rebuffer5670 (.A(net5981),
    .Y(net5670));
 BUFx3_ASAP7_75t_R rebuffer5671 (.A(_03720_),
    .Y(net5671));
 BUFx3_ASAP7_75t_R rebuffer5672 (.A(_03736_),
    .Y(net5672));
 BUFx3_ASAP7_75t_R rebuffer5673 (.A(_03354_),
    .Y(net5673));
 BUFx3_ASAP7_75t_R rebuffer5674 (.A(_03610_),
    .Y(net5674));
 BUFx6f_ASAP7_75t_R rebuffer5675 (.A(_03610_),
    .Y(net5675));
 BUFx3_ASAP7_75t_R rebuffer5676 (.A(_03691_),
    .Y(net5676));
 BUFx3_ASAP7_75t_R rebuffer5677 (.A(_03900_),
    .Y(net5677));
 BUFx6f_ASAP7_75t_R rebuffer5678 (.A(_03728_),
    .Y(net5678));
 BUFx3_ASAP7_75t_R rebuffer5679 (.A(_03601_),
    .Y(net5679));
 BUFx3_ASAP7_75t_R rebuffer5680 (.A(_03354_),
    .Y(net5680));
 BUFx3_ASAP7_75t_R rebuffer5681 (.A(_03833_),
    .Y(net5681));
 BUFx3_ASAP7_75t_R rebuffer5682 (.A(_03727_),
    .Y(net5682));
 BUFx3_ASAP7_75t_R rebuffer5683 (.A(net5695),
    .Y(net5683));
 BUFx3_ASAP7_75t_R rebuffer5684 (.A(_04025_),
    .Y(net5684));
 BUFx3_ASAP7_75t_R rebuffer5685 (.A(_04055_),
    .Y(net5685));
 BUFx6f_ASAP7_75t_R rebuffer5686 (.A(_03737_),
    .Y(net5686));
 BUFx3_ASAP7_75t_R rebuffer5687 (.A(_04043_),
    .Y(net5687));
 BUFx3_ASAP7_75t_R rebuffer5688 (.A(_04054_),
    .Y(net5688));
 BUFx3_ASAP7_75t_R rebuffer5689 (.A(_03541_),
    .Y(net5689));
 BUFx3_ASAP7_75t_R rebuffer5690 (.A(_03557_),
    .Y(net5690));
 BUFx3_ASAP7_75t_R rebuffer5691 (.A(_03602_),
    .Y(net5691));
 BUFx3_ASAP7_75t_R rebuffer5692 (.A(_02495_),
    .Y(net5692));
 BUFx3_ASAP7_75t_R rebuffer5693 (.A(_04108_),
    .Y(net5693));
 BUFx3_ASAP7_75t_R rebuffer5694 (.A(_03746_),
    .Y(net5694));
 BUFx3_ASAP7_75t_R rebuffer5695 (.A(_03385_),
    .Y(net5695));
 BUFx3_ASAP7_75t_R rebuffer5696 (.A(_03385_),
    .Y(net5696));
 BUFx6f_ASAP7_75t_R rebuffer5697 (.A(_03378_),
    .Y(net5697));
 BUFx3_ASAP7_75t_R rebuffer5698 (.A(_03493_),
    .Y(net5698));
 BUFx3_ASAP7_75t_R rebuffer5699 (.A(_03498_),
    .Y(net5699));
 BUFx3_ASAP7_75t_R rebuffer5700 (.A(_03717_),
    .Y(net5700));
 BUFx3_ASAP7_75t_R rebuffer5701 (.A(_03649_),
    .Y(net5701));
 BUFx3_ASAP7_75t_R rebuffer5702 (.A(_04096_),
    .Y(net5702));
 BUFx3_ASAP7_75t_R rebuffer5703 (.A(_03751_),
    .Y(net5703));
 BUFx3_ASAP7_75t_R rebuffer5704 (.A(_03644_),
    .Y(net5704));
 BUFx3_ASAP7_75t_R rebuffer5705 (.A(_03574_),
    .Y(net5705));
 BUFx3_ASAP7_75t_R rebuffer5706 (.A(_03444_),
    .Y(net5706));
 BUFx3_ASAP7_75t_R rebuffer5707 (.A(_03241_),
    .Y(net5707));
 BUFx3_ASAP7_75t_R rebuffer5708 (.A(net4965),
    .Y(net5708));
 BUFx3_ASAP7_75t_R rebuffer5709 (.A(net5708),
    .Y(net5709));
 BUFx3_ASAP7_75t_R rebuffer5710 (.A(_00533_),
    .Y(net5710));
 BUFx3_ASAP7_75t_R rebuffer5714 (.A(_03225_),
    .Y(net5714));
 BUFx3_ASAP7_75t_R rebuffer5715 (.A(_04074_),
    .Y(net5715));
 BUFx3_ASAP7_75t_R rebuffer5716 (.A(_03299_),
    .Y(net5716));
 BUFx3_ASAP7_75t_R rebuffer5718 (.A(net6011),
    .Y(net5718));
 BUFx3_ASAP7_75t_R rebuffer5719 (.A(_04086_),
    .Y(net5719));
 BUFx3_ASAP7_75t_R rebuffer5720 (.A(_04091_),
    .Y(net5720));
 BUFx3_ASAP7_75t_R rebuffer5728 (.A(_04140_),
    .Y(net5728));
 BUFx3_ASAP7_75t_R rebuffer5757 (.A(_01716_),
    .Y(net5757));
 BUFx3_ASAP7_75t_R rebuffer5758 (.A(_01058_),
    .Y(net5758));
 BUFx3_ASAP7_75t_R rebuffer5759 (.A(_02340_),
    .Y(net5759));
 BUFx3_ASAP7_75t_R rebuffer5760 (.A(_01878_),
    .Y(net5760));
 BUFx3_ASAP7_75t_R rebuffer5761 (.A(_00078_),
    .Y(net5761));
 BUFx6f_ASAP7_75t_R rebuffer5762 (.A(_01739_),
    .Y(net5762));
 BUFx3_ASAP7_75t_R rebuffer5763 (.A(_01705_),
    .Y(net5763));
 BUFx3_ASAP7_75t_R rebuffer5764 (.A(_01739_),
    .Y(net5764));
 BUFx6f_ASAP7_75t_R rebuffer5765 (.A(_02053_),
    .Y(net5765));
 BUFx3_ASAP7_75t_R rebuffer5766 (.A(_01674_),
    .Y(net5766));
 BUFx3_ASAP7_75t_R rebuffer5767 (.A(_01230_),
    .Y(net5767));
 BUFx3_ASAP7_75t_R rebuffer5768 (.A(_01666_),
    .Y(net5768));
 BUFx3_ASAP7_75t_R rebuffer5769 (.A(_02327_),
    .Y(net5769));
 BUFx3_ASAP7_75t_R rebuffer5770 (.A(_01941_),
    .Y(net5770));
 BUFx3_ASAP7_75t_R rebuffer5771 (.A(_01693_),
    .Y(net5771));
 BUFx3_ASAP7_75t_R rebuffer5772 (.A(_00524_),
    .Y(net5772));
 BUFx3_ASAP7_75t_R rebuffer5773 (.A(_01993_),
    .Y(net5773));
 BUFx3_ASAP7_75t_R rebuffer5787 (.A(_01831_),
    .Y(net5787));
 BUFx3_ASAP7_75t_R rebuffer5819 (.A(net3416),
    .Y(net5819));
 BUFx3_ASAP7_75t_R rebuffer5820 (.A(net3416),
    .Y(net5820));
 BUFx3_ASAP7_75t_R rebuffer5821 (.A(_02326_),
    .Y(net5821));
 BUFx3_ASAP7_75t_R rebuffer5822 (.A(net3539),
    .Y(net5822));
 BUFx3_ASAP7_75t_R rebuffer5876 (.A(_02343_),
    .Y(net5876));
 BUFx3_ASAP7_75t_R rebuffer5877 (.A(_02343_),
    .Y(net5877));
 BUFx3_ASAP7_75t_R rebuffer5887 (.A(_02250_),
    .Y(net5887));
 BUFx3_ASAP7_75t_R rebuffer5888 (.A(_01687_),
    .Y(net5888));
 BUFx3_ASAP7_75t_R rebuffer5889 (.A(net3805),
    .Y(net5889));
 BUFx3_ASAP7_75t_R rebuffer5894 (.A(_02230_),
    .Y(net5894));
 BUFx12f_ASAP7_75t_R clone5895 (.A(net5372),
    .Y(net5895));
 BUFx3_ASAP7_75t_R rebuffer5902 (.A(_02351_),
    .Y(net5902));
 BUFx6f_ASAP7_75t_R rebuffer5903 (.A(net5419),
    .Y(net5903));
 BUFx12f_ASAP7_75t_R clone5912 (.A(_04330_),
    .Y(net5912));
 BUFx3_ASAP7_75t_R rebuffer5913 (.A(_01454_),
    .Y(net5913));
 BUFx3_ASAP7_75t_R rebuffer5914 (.A(\u_window_buffer.internal_read_ptr[2] ),
    .Y(net5914));
 BUFx3_ASAP7_75t_R rebuffer5917 (.A(_01425_),
    .Y(net5917));
 BUFx3_ASAP7_75t_R rebuffer5918 (.A(_01450_),
    .Y(net5918));
 BUFx12f_ASAP7_75t_R clone5920 (.A(_04330_),
    .Y(net5920));
 BUFx6f_ASAP7_75t_R rebuffer5923 (.A(net2699),
    .Y(net5923));
 BUFx3_ASAP7_75t_R rebuffer5924 (.A(_06216_),
    .Y(net5924));
 BUFx3_ASAP7_75t_R rebuffer5933 (.A(_05869_),
    .Y(net5933));
 BUFx3_ASAP7_75t_R rebuffer5934 (.A(_05991_),
    .Y(net5934));
 BUFx3_ASAP7_75t_R rebuffer5935 (.A(_05902_),
    .Y(net5935));
 BUFx3_ASAP7_75t_R rebuffer5936 (.A(_06137_),
    .Y(net5936));
 BUFx3_ASAP7_75t_R rebuffer5937 (.A(_05893_),
    .Y(net5937));
 BUFx3_ASAP7_75t_R rebuffer5938 (.A(_05677_),
    .Y(net5938));
 BUFx3_ASAP7_75t_R rebuffer5939 (.A(_05827_),
    .Y(net5939));
 BUFx3_ASAP7_75t_R rebuffer5940 (.A(_05995_),
    .Y(net5940));
 BUFx3_ASAP7_75t_R rebuffer5941 (.A(_05966_),
    .Y(net5941));
 BUFx3_ASAP7_75t_R rebuffer5957 (.A(_06448_),
    .Y(net5957));
 BUFx3_ASAP7_75t_R rebuffer5958 (.A(_06350_),
    .Y(net5958));
 BUFx3_ASAP7_75t_R rebuffer5959 (.A(_05649_),
    .Y(net5959));
 BUFx3_ASAP7_75t_R rebuffer5960 (.A(_05540_),
    .Y(net5960));
 BUFx3_ASAP7_75t_R rebuffer5961 (.A(_05785_),
    .Y(net5961));
 BUFx3_ASAP7_75t_R rebuffer5964 (.A(_06411_),
    .Y(net5964));
 BUFx3_ASAP7_75t_R rebuffer5972 (.A(_03860_),
    .Y(net5972));
 BUFx3_ASAP7_75t_R rebuffer5973 (.A(_03562_),
    .Y(net5973));
 BUFx6f_ASAP7_75t_R rebuffer5974 (.A(_03598_),
    .Y(net5974));
 BUFx3_ASAP7_75t_R rebuffer5975 (.A(_03439_),
    .Y(net5975));
 BUFx3_ASAP7_75t_R rebuffer5976 (.A(_04038_),
    .Y(net5976));
 BUFx3_ASAP7_75t_R rebuffer5977 (.A(_03358_),
    .Y(net5977));
 BUFx3_ASAP7_75t_R rebuffer5978 (.A(_03651_),
    .Y(net5978));
 BUFx3_ASAP7_75t_R rebuffer5979 (.A(_03470_),
    .Y(net5979));
 BUFx3_ASAP7_75t_R rebuffer5980 (.A(_03779_),
    .Y(net5980));
 BUFx6f_ASAP7_75t_R rebuffer5981 (.A(_03764_),
    .Y(net5981));
 BUFx3_ASAP7_75t_R rebuffer5982 (.A(_03663_),
    .Y(net5982));
 BUFx3_ASAP7_75t_R rebuffer5983 (.A(_04121_),
    .Y(net5983));
 BUFx3_ASAP7_75t_R rebuffer5984 (.A(_03602_),
    .Y(net5984));
 BUFx3_ASAP7_75t_R rebuffer5985 (.A(_03565_),
    .Y(net5985));
 BUFx3_ASAP7_75t_R rebuffer5986 (.A(_03597_),
    .Y(net5986));
 BUFx3_ASAP7_75t_R rebuffer5987 (.A(_03438_),
    .Y(net5987));
 BUFx3_ASAP7_75t_R rebuffer5988 (.A(_03685_),
    .Y(net5988));
 BUFx3_ASAP7_75t_R rebuffer5996 (.A(_03651_),
    .Y(net5996));
 BUFx3_ASAP7_75t_R rebuffer5997 (.A(_03615_),
    .Y(net5997));
 BUFx3_ASAP7_75t_R rebuffer5998 (.A(_03790_),
    .Y(net5998));
 BUFx3_ASAP7_75t_R rebuffer5999 (.A(_03636_),
    .Y(net5999));
 BUFx3_ASAP7_75t_R rebuffer6000 (.A(_03408_),
    .Y(net6000));
 BUFx3_ASAP7_75t_R rebuffer6003 (.A(net3314),
    .Y(net6003));
 BUFx3_ASAP7_75t_R rebuffer6010 (.A(_03452_),
    .Y(net6010));
 BUFx3_ASAP7_75t_R rebuffer6011 (.A(_04078_),
    .Y(net6011));
 BUFx3_ASAP7_75t_R rebuffer6030 (.A(_02818_),
    .Y(net6030));
 BUFx3_ASAP7_75t_R rebuffer6033 (.A(net6037),
    .Y(net6033));
 BUFx3_ASAP7_75t_R rebuffer6034 (.A(net6037),
    .Y(net6034));
 BUFx6f_ASAP7_75t_R rebuffer6035 (.A(net3998),
    .Y(net6035));
 BUFx3_ASAP7_75t_R rebuffer6036 (.A(net6037),
    .Y(net6036));
 BUFx6f_ASAP7_75t_R clone6037 (.A(net6040),
    .Y(net6037));
 BUFx3_ASAP7_75t_R rebuffer6038 (.A(_02896_),
    .Y(net6038));
 BUFx3_ASAP7_75t_R rebuffer6039 (.A(net4018),
    .Y(net6039));
 BUFx3_ASAP7_75t_R rebuffer6040 (.A(_02899_),
    .Y(net6040));
 BUFx3_ASAP7_75t_R rebuffer6041 (.A(_02812_),
    .Y(net6041));
 BUFx3_ASAP7_75t_R rebuffer6042 (.A(_02804_),
    .Y(net6042));
 BUFx3_ASAP7_75t_R rebuffer6043 (.A(net3999),
    .Y(net6043));
endmodule
