module DCT (
    ports
);

logic signed [15:0] cos_table [40][12] = '{
    '{ 16'sd32767, 16'sd32742, 16'sd32666, 16'sd32540, 16'sd32364, 16'sd32138, 16'sd31862, 16'sd31537, 16'sd31164, 16'sd30742, 16'sd30273, 16'sd29758 },
    '{ 16'sd32767, 16'sd32540, 16'sd31862, 16'sd30742, 16'sd29196, 16'sd27245, 16'sd24916, 16'sd22242, 16'sd19260, 16'sd16011, 16'sd12539, 16'sd8894 },
    '{ 16'sd32767, 16'sd32138, 16'sd30273, 16'sd27245, 16'sd23170, 16'sd18204, 16'sd12539, 16'sd6392, 16'sd0, 16'sd-6392, 16'sd-12539, 16'sd-18204 },
    '{ 16'sd32767, 16'sd31537, 16'sd27939, 16'sd22242, 16'sd14876, 16'sd6392, 16'sd-2570, 16'sd-11341, 16'sd-19260, 16'sd-25733, 16'sd-30273, 16'sd-32540 },
    '{ 16'sd32767, 16'sd30742, 16'sd24916, 16'sd16011, 16'sd5126, 16'sd-6392, 16'sd-17121, 16'sd-25733, 16'sd-31164, 16'sd-32742, 16'sd-30273, 16'sd-24062 },
    '{ 16'sd32767, 16'sd29758, 16'sd21281, 16'sd8894, 16'sd-5126, 16'sd-18204, 16'sd-27939, 16'sd-32540, 16'sd-31164, 16'sd-24062, 16'sd-12539, 16'sd1286 },
    '{ 16'sd32767, 16'sd28589, 16'sd17121, 16'sd1286, 16'sd-14876, 16'sd-27245, 16'sd-32666, 16'sd-29758, 16'sd-19260, 16'sd-3851, 16'sd12539, 16'sd25733 },
    '{ 16'sd32767, 16'sd27245, 16'sd12539, 16'sd-6392, 16'sd-23170, 16'sd-32138, 16'sd-30273, 16'sd-18204, 16'sd0, 16'sd18204, 16'sd30273, 16'sd32138 },
    '{ 16'sd32767, 16'sd25733, 16'sd7649, 16'sd-13718, 16'sd-29196, 16'sd-32138, 16'sd-21281, 16'sd-1286, 16'sd19260, 16'sd31537, 16'sd30273, 16'sd16011 },
    '{ 16'sd32767, 16'sd24062, 16'sd2570, 16'sd-20286, 16'sd-32364, 16'sd-27245, 16'sd-7649, 16'sd16011, 16'sd31164, 16'sd29758, 16'sd12539, 16'sd-11341 },
    '{ 16'sd32767, 16'sd22242, 16'sd-2570, 16'sd-25733, 16'sd-32364, 16'sd-18204, 16'sd7649, 16'sd28589, 16'sd31164, 16'sd13718, 16'sd-12539, 16'sd-30742 },
    '{ 16'sd32767, 16'sd20286, 16'sd-7649, 16'sd-29758, 16'sd-29196, 16'sd-6392, 16'sd21281, 16'sd32742, 16'sd19260, 16'sd-8894, 16'sd-30273, 16'sd-28589 },
    '{ 16'sd32767, 16'sd18204, 16'sd-12539, 16'sd-32138, 16'sd-23170, 16'sd6392, 16'sd30273, 16'sd27245, 16'sd0, 16'sd-27245, 16'sd-30273, 16'sd-6392 },
    '{ 16'sd32767, 16'sd16011, 16'sd-17121, 16'sd-32742, 16'sd-14876, 16'sd18204, 16'sd32666, 16'sd13718, 16'sd-19260, 16'sd-32540, 16'sd-12539, 16'sd20286 },
    '{ 16'sd32767, 16'sd13718, 16'sd-21281, 16'sd-31537, 16'sd-5126, 16'sd27245, 16'sd27939, 16'sd-3851, 16'sd-31164, 16'sd-22242, 16'sd12539, 16'sd32742 },
    '{ 16'sd32767, 16'sd11341, 16'sd-24916, 16'sd-28589, 16'sd5126, 16'sd32138, 16'sd17121, 16'sd-20286, 16'sd-31164, 16'sd-1286, 16'sd30273, 16'sd22242 },
    '{ 16'sd32767, 16'sd8894, 16'sd-27939, 16'sd-24062, 16'sd14876, 16'sd32138, 16'sd2570, 16'sd-30742, 16'sd-19260, 16'sd20286, 16'sd30273, 16'sd-3851 },
    '{ 16'sd32767, 16'sd6392, 16'sd-30273, 16'sd-18204, 16'sd23170, 16'sd27245, 16'sd-12539, 16'sd-32138, 16'sd0, 16'sd32138, 16'sd12539, 16'sd-27245 },
    '{ 16'sd32767, 16'sd3851, 16'sd-31862, 16'sd-11341, 16'sd29196, 16'sd18204, 16'sd-24916, 16'sd-24062, 16'sd19260, 16'sd28589, 16'sd-12539, 16'sd-31537 },
    '{ 16'sd32767, 16'sd1286, 16'sd-32666, 16'sd-3851, 16'sd32364, 16'sd6392, 16'sd-31862, 16'sd-8894, 16'sd31164, 16'sd11341, 16'sd-30273, 16'sd-13718 },
    '{ 16'sd32767, 16'sd-1286, 16'sd-32666, 16'sd3851, 16'sd32364, 16'sd-6392, 16'sd-31862, 16'sd8894, 16'sd31164, 16'sd-11341, 16'sd-30273, 16'sd13718 },
    '{ 16'sd32767, 16'sd-3851, 16'sd-31862, 16'sd11341, 16'sd29196, 16'sd-18204, 16'sd-24916, 16'sd24062, 16'sd19260, 16'sd-28589, 16'sd-12539, 16'sd31537 },
    '{ 16'sd32767, 16'sd-6392, 16'sd-30273, 16'sd18204, 16'sd23170, 16'sd-27245, 16'sd-12539, 16'sd32138, 16'sd0, 16'sd-32138, 16'sd12539, 16'sd27245 },
    '{ 16'sd32767, 16'sd-8894, 16'sd-27939, 16'sd24062, 16'sd14876, 16'sd-32138, 16'sd2570, 16'sd30742, 16'sd-19260, 16'sd-20286, 16'sd30273, 16'sd3851 },
    '{ 16'sd32767, 16'sd-11341, 16'sd-24916, 16'sd28589, 16'sd5126, 16'sd-32138, 16'sd17121, 16'sd20286, 16'sd-31164, 16'sd1286, 16'sd30273, 16'sd-22242 },
    '{ 16'sd32767, 16'sd-13718, 16'sd-21281, 16'sd31537, 16'sd-5126, 16'sd-27245, 16'sd27939, 16'sd3851, 16'sd-31164, 16'sd22242, 16'sd12539, 16'sd-32742 },
    '{ 16'sd32767, 16'sd-16011, 16'sd-17121, 16'sd32742, 16'sd-14876, 16'sd-18204, 16'sd32666, 16'sd-13718, 16'sd-19260, 16'sd32540, 16'sd-12539, 16'sd-20286 },
    '{ 16'sd32767, 16'sd-18204, 16'sd-12539, 16'sd32138, 16'sd-23170, 16'sd-6392, 16'sd30273, 16'sd-27245, 16'sd0, 16'sd27245, 16'sd-30273, 16'sd6392 },
    '{ 16'sd32767, 16'sd-20286, 16'sd-7649, 16'sd29758, 16'sd-29196, 16'sd6392, 16'sd21281, 16'sd-32742, 16'sd19260, 16'sd8894, 16'sd-30273, 16'sd28589 },
    '{ 16'sd32767, 16'sd-22242, 16'sd-2570, 16'sd25733, 16'sd-32364, 16'sd18204, 16'sd7649, 16'sd-28589, 16'sd31164, 16'sd-13718, 16'sd-12539, 16'sd30742 },
    '{ 16'sd32767, 16'sd-24062, 16'sd2570, 16'sd20286, 16'sd-32364, 16'sd27245, 16'sd-7649, 16'sd-16011, 16'sd31164, 16'sd-29758, 16'sd12539, 16'sd11341 },
    '{ 16'sd32767, 16'sd-25733, 16'sd7649, 16'sd13718, 16'sd-29196, 16'sd32138, 16'sd-21281, 16'sd1286, 16'sd19260, 16'sd-31537, 16'sd30273, 16'sd-16011 },
    '{ 16'sd32767, 16'sd-27245, 16'sd12539, 16'sd6392, 16'sd-23170, 16'sd32138, 16'sd-30273, 16'sd18204, 16'sd0, 16'sd-18204, 16'sd30273, 16'sd-32138 },
    '{ 16'sd32767, 16'sd-28589, 16'sd17121, 16'sd-1286, 16'sd-14876, 16'sd27245, 16'sd-32666, 16'sd29758, 16'sd-19260, 16'sd3851, 16'sd12539, 16'sd-25733 },
    '{ 16'sd32767, 16'sd-29758, 16'sd21281, 16'sd-8894, 16'sd-5126, 16'sd18204, 16'sd-27939, 16'sd32540, 16'sd-31164, 16'sd24062, 16'sd-12539, 16'sd-1286 },
    '{ 16'sd32767, 16'sd-30742, 16'sd24916, 16'sd-16011, 16'sd5126, 16'sd6392, 16'sd-17121, 16'sd25733, 16'sd-31164, 16'sd32742, 16'sd-30273, 16'sd24062 },
    '{ 16'sd32767, 16'sd-31537, 16'sd27939, 16'sd-22242, 16'sd14876, 16'sd-6392, 16'sd-2570, 16'sd11341, 16'sd-19260, 16'sd25733, 16'sd-30273, 16'sd32540 },
    '{ 16'sd32767, 16'sd-32138, 16'sd30273, 16'sd-27245, 16'sd23170, 16'sd-18204, 16'sd12539, 16'sd-6392, 16'sd0, 16'sd6392, 16'sd-12539, 16'sd18204 },
    '{ 16'sd32767, 16'sd-32540, 16'sd31862, 16'sd-30742, 16'sd29196, 16'sd-27245, 16'sd24916, 16'sd-22242, 16'sd19260, 16'sd-16011, 16'sd12539, 16'sd-8894 },
    '{ 16'sd32767, 16'sd-32742, 16'sd32666, 16'sd-32540, 16'sd32364, 16'sd-32138, 16'sd31862, 16'sd-31537, 16'sd31164, 16'sd-30742, 16'sd30273, 16'sd-29758 }
};
    
endmodule