`timescale 1ns/1ps

module MEL #(
    parameter NUM_FILTERS = 40
) (
    input  logic clk,
    input  logic rst_n,
);
    
endmodule